VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt08-ssp-opamp
  CLASS BLOCK ;
  FOREIGN tt08-ssp-opamp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.280900 ;
    PORT
      LAYER li1 ;
        RECT 131.060 67.090 131.485 67.285 ;
        RECT 131.060 66.880 131.490 67.090 ;
        RECT 131.060 66.655 131.485 66.880 ;
        RECT 131.220 65.345 131.485 66.655 ;
        RECT 130.830 65.075 131.485 65.345 ;
      LAYER met1 ;
        RECT 132.960 67.120 152.750 67.790 ;
        RECT 131.150 66.880 152.750 67.120 ;
        RECT 131.150 66.850 131.550 66.880 ;
        RECT 132.960 66.800 152.750 66.880 ;
        RECT 150.790 66.710 152.750 66.800 ;
      LAYER met2 ;
        RECT 150.840 66.660 152.700 67.840 ;
      LAYER met3 ;
        RECT 150.790 66.685 152.750 67.815 ;
      LAYER met4 ;
        RECT 150.835 67.710 152.705 67.795 ;
        RECT 150.835 66.705 152.710 67.710 ;
        RECT 151.810 0.000 152.710 66.705 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.750000 ;
    ANTENNADIFFAREA 18.039999 ;
    PORT
      LAYER li1 ;
        RECT 126.770 89.320 126.940 89.650 ;
        RECT 136.320 88.840 136.560 89.180 ;
        RECT 126.770 88.360 126.940 88.690 ;
        RECT 136.320 87.880 136.490 88.210 ;
        RECT 113.450 84.280 113.780 84.450 ;
        RECT 114.410 84.280 114.740 84.450 ;
        RECT 123.620 77.865 123.790 79.905 ;
        RECT 124.580 77.865 124.750 79.905 ;
        RECT 125.540 77.865 125.710 79.905 ;
        RECT 112.970 74.640 113.300 74.810 ;
        RECT 113.930 74.640 114.260 74.810 ;
        RECT 121.000 70.165 121.170 71.205 ;
        RECT 114.850 69.450 115.150 69.490 ;
        RECT 114.840 69.280 115.170 69.450 ;
        RECT 114.850 69.250 115.150 69.280 ;
        RECT 117.570 68.490 117.900 68.660 ;
        RECT 118.530 68.490 118.860 68.660 ;
        RECT 102.840 58.735 103.010 66.775 ;
        RECT 103.800 58.735 103.970 66.775 ;
        RECT 104.760 58.735 104.930 66.775 ;
        RECT 105.720 58.735 105.890 66.775 ;
        RECT 106.680 58.735 106.850 66.775 ;
        RECT 107.640 58.735 107.810 66.775 ;
        RECT 117.090 65.940 117.420 66.110 ;
        RECT 118.050 65.940 118.380 66.110 ;
        RECT 119.010 65.940 119.340 66.110 ;
        RECT 114.840 65.640 115.170 65.810 ;
        RECT 104.590 54.680 104.760 55.720 ;
      LAYER met1 ;
        RECT 116.170 91.020 117.460 91.130 ;
        RECT 116.095 91.010 136.600 91.020 ;
        RECT 116.095 90.410 136.610 91.010 ;
        RECT 112.820 84.750 115.370 84.830 ;
        RECT 116.170 84.750 117.460 90.410 ;
        RECT 126.650 89.650 126.970 90.410 ;
        RECT 126.650 88.370 126.980 89.650 ;
        RECT 136.340 89.170 136.610 90.410 ;
        RECT 126.660 88.360 126.980 88.370 ;
        RECT 136.290 87.880 136.610 89.170 ;
        RECT 136.290 87.870 136.570 87.880 ;
        RECT 112.820 84.320 117.460 84.750 ;
        RECT 112.820 84.290 117.050 84.320 ;
        RECT 112.820 84.190 115.370 84.290 ;
        RECT 112.280 74.870 114.830 74.880 ;
        RECT 116.090 74.870 116.490 84.290 ;
        RECT 123.590 79.700 123.820 79.885 ;
        RECT 123.450 79.180 123.920 79.700 ;
        RECT 124.550 79.670 124.780 79.885 ;
        RECT 123.590 77.885 123.820 79.180 ;
        RECT 124.490 79.150 124.860 79.670 ;
        RECT 125.510 79.660 125.740 79.885 ;
        RECT 124.550 77.885 124.780 79.150 ;
        RECT 125.420 79.140 125.790 79.660 ;
        RECT 125.510 77.885 125.740 79.140 ;
        RECT 112.280 74.440 118.040 74.870 ;
        RECT 112.280 74.240 114.830 74.440 ;
        RECT 112.630 69.720 113.900 74.240 ;
        RECT 120.840 70.150 121.250 71.200 ;
        RECT 112.600 69.690 117.660 69.720 ;
        RECT 112.550 69.190 117.660 69.690 ;
        RECT 112.550 68.990 113.820 69.190 ;
        RECT 112.550 68.380 113.900 68.990 ;
        RECT 117.120 68.800 117.630 69.190 ;
        RECT 117.120 68.460 120.270 68.800 ;
        RECT 117.150 68.440 120.270 68.460 ;
        RECT 112.630 67.140 113.900 68.380 ;
        RECT 102.810 66.740 103.040 66.755 ;
        RECT 102.720 64.460 103.110 66.740 ;
        RECT 103.770 66.720 104.000 66.755 ;
        RECT 104.730 66.750 104.960 66.755 ;
        RECT 102.810 58.755 103.040 64.460 ;
        RECT 103.680 64.440 104.070 66.720 ;
        RECT 104.650 64.470 105.040 66.750 ;
        RECT 105.690 66.740 105.920 66.755 ;
        RECT 106.650 66.740 106.880 66.755 ;
        RECT 103.770 58.755 104.000 64.440 ;
        RECT 104.730 58.755 104.960 64.470 ;
        RECT 105.610 64.460 106.000 66.740 ;
        RECT 106.580 64.460 106.970 66.740 ;
        RECT 107.610 66.720 107.840 66.755 ;
        RECT 105.690 58.755 105.920 64.460 ;
        RECT 106.650 58.755 106.880 64.460 ;
        RECT 107.540 64.440 107.930 66.720 ;
        RECT 112.630 65.910 113.890 67.140 ;
        RECT 119.820 66.150 120.270 68.440 ;
        RECT 112.600 65.890 114.590 65.910 ;
        RECT 112.600 65.870 116.000 65.890 ;
        RECT 116.670 65.870 120.270 66.150 ;
        RECT 112.600 65.850 120.270 65.870 ;
        RECT 112.600 65.830 120.250 65.850 ;
        RECT 112.600 65.590 117.000 65.830 ;
        RECT 118.640 65.820 119.710 65.830 ;
        RECT 112.600 65.540 116.830 65.590 ;
        RECT 112.600 65.530 116.000 65.540 ;
        RECT 114.010 65.510 116.000 65.530 ;
        RECT 107.610 58.755 107.840 64.440 ;
        RECT 104.560 55.040 104.790 55.700 ;
        RECT 104.390 54.760 104.790 55.040 ;
        RECT 104.560 54.700 104.790 54.760 ;
      LAYER met2 ;
        RECT 123.370 79.750 123.740 79.850 ;
        RECT 123.370 79.720 123.870 79.750 ;
        RECT 123.370 79.180 125.790 79.720 ;
        RECT 123.370 79.130 123.870 79.180 ;
        RECT 120.850 73.730 121.260 73.780 ;
        RECT 123.370 73.730 123.740 79.130 ;
        RECT 124.540 79.100 124.810 79.180 ;
        RECT 125.470 79.090 125.740 79.180 ;
        RECT 120.800 73.100 124.070 73.730 ;
        RECT 120.850 71.160 121.260 73.100 ;
        RECT 112.670 70.250 121.260 71.160 ;
        RECT 112.670 70.120 121.240 70.250 ;
        RECT 112.710 69.760 113.640 70.120 ;
        RECT 120.890 70.100 121.200 70.120 ;
        RECT 112.710 69.390 113.630 69.760 ;
        RECT 112.650 68.120 113.630 69.390 ;
        RECT 110.180 67.760 110.790 67.990 ;
        RECT 112.710 67.830 113.630 68.120 ;
        RECT 112.680 67.760 113.630 67.830 ;
        RECT 110.180 66.860 113.690 67.760 ;
        RECT 102.770 66.630 103.060 66.790 ;
        RECT 103.730 66.630 104.020 66.770 ;
        RECT 104.700 66.630 104.990 66.800 ;
        RECT 105.660 66.630 105.950 66.790 ;
        RECT 106.630 66.630 106.920 66.790 ;
        RECT 107.590 66.630 107.880 66.770 ;
        RECT 102.620 65.410 107.930 66.630 ;
        RECT 110.180 65.560 110.790 66.860 ;
        RECT 112.680 66.810 113.630 66.860 ;
        RECT 112.680 66.660 113.590 66.810 ;
        RECT 110.180 65.410 110.780 65.560 ;
        RECT 102.620 64.760 110.790 65.410 ;
        RECT 102.620 64.470 107.930 64.760 ;
        RECT 102.770 64.410 103.060 64.470 ;
        RECT 103.730 64.390 104.020 64.470 ;
        RECT 104.700 64.420 104.990 64.470 ;
        RECT 105.660 64.410 105.950 64.470 ;
        RECT 106.630 64.410 106.920 64.470 ;
        RECT 107.590 64.390 107.880 64.470 ;
        RECT 110.180 56.270 110.780 64.760 ;
        RECT 110.180 55.140 110.900 56.270 ;
        RECT 104.420 54.730 110.900 55.140 ;
        RECT 104.420 54.700 110.860 54.730 ;
      LAYER met3 ;
        RECT 112.600 68.145 113.620 69.365 ;
        RECT 115.690 45.260 117.120 46.470 ;
        RECT 115.790 3.740 116.690 45.260 ;
        RECT 131.310 3.740 133.500 3.830 ;
        RECT 115.790 2.840 133.500 3.740 ;
        RECT 131.310 2.830 133.500 2.840 ;
      LAYER met4 ;
        RECT 112.645 69.130 113.575 69.345 ;
        RECT 116.250 69.130 117.030 69.190 ;
        RECT 112.610 68.160 117.030 69.130 ;
        RECT 116.250 46.475 117.030 68.160 ;
        RECT 115.735 45.255 117.075 46.475 ;
        RECT 131.355 2.825 133.455 3.835 ;
        RECT 132.490 0.000 133.390 2.825 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.751700 ;
    PORT
      LAYER li1 ;
        RECT 106.400 21.020 106.570 26.060 ;
        RECT 107.980 21.020 108.150 26.060 ;
        RECT 109.560 21.020 109.730 26.060 ;
        RECT 105.440 12.210 105.610 16.160 ;
        RECT 107.020 12.210 107.190 16.160 ;
        RECT 108.600 12.210 108.770 16.160 ;
      LAYER met1 ;
        RECT 106.370 24.910 106.600 26.040 ;
        RECT 107.950 24.910 108.180 26.040 ;
        RECT 109.530 24.910 109.760 26.040 ;
        RECT 106.370 24.760 106.700 24.910 ;
        RECT 106.370 22.750 106.810 24.760 ;
        RECT 106.370 21.040 106.600 22.750 ;
        RECT 107.950 22.690 108.270 24.910 ;
        RECT 109.530 22.690 109.850 24.910 ;
        RECT 107.950 21.040 108.180 22.690 ;
        RECT 109.530 21.040 109.760 22.690 ;
        RECT 105.410 15.520 105.640 16.140 ;
        RECT 106.990 15.540 107.220 16.140 ;
        RECT 108.570 15.550 108.800 16.140 ;
        RECT 105.410 13.300 105.810 15.520 ;
        RECT 106.990 13.320 107.400 15.540 ;
        RECT 108.570 13.330 108.980 15.550 ;
        RECT 105.410 12.230 105.640 13.300 ;
        RECT 106.990 12.230 107.220 13.320 ;
        RECT 108.570 12.230 108.800 13.330 ;
      LAYER met2 ;
        RECT 106.120 22.990 109.910 24.910 ;
        RECT 106.120 22.690 114.850 22.990 ;
        RECT 106.750 21.390 114.850 22.690 ;
        RECT 106.780 15.630 108.430 21.390 ;
        RECT 105.070 13.160 109.210 15.630 ;
      LAYER met3 ;
        RECT 112.300 21.390 114.850 22.990 ;
      LAYER met4 ;
        RECT 118.245 22.990 147.855 43.895 ;
        RECT 112.300 21.390 147.855 22.990 ;
        RECT 113.170 0.000 114.070 21.390 ;
        RECT 118.245 14.285 147.855 21.390 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 16.820000 ;
    PORT
      LAYER li1 ;
        RECT 33.680 9.880 33.850 19.920 ;
        RECT 36.260 9.880 36.430 19.920 ;
        RECT 41.110 18.535 41.280 37.575 ;
        RECT 42.090 18.535 42.260 37.575 ;
      LAYER met1 ;
        RECT 33.650 19.490 33.880 19.900 ;
        RECT 33.450 18.750 34.110 19.490 ;
        RECT 36.230 19.430 36.460 19.900 ;
        RECT 41.080 19.500 41.310 37.555 ;
        RECT 42.060 19.510 42.290 37.555 ;
        RECT 33.650 9.900 33.880 18.750 ;
        RECT 36.030 18.690 36.690 19.430 ;
        RECT 40.980 18.750 41.410 19.500 ;
        RECT 41.960 18.760 42.390 19.510 ;
        RECT 36.230 9.900 36.460 18.690 ;
        RECT 41.080 18.555 41.310 18.750 ;
        RECT 42.060 18.555 42.290 18.760 ;
        RECT 84.280 17.290 92.610 21.970 ;
      LAYER met2 ;
        RECT 84.330 20.340 92.560 22.020 ;
        RECT 78.490 20.190 92.560 20.340 ;
        RECT 33.390 20.180 39.800 20.190 ;
        RECT 40.610 20.180 92.560 20.190 ;
        RECT 33.390 18.520 92.560 20.180 ;
        RECT 33.390 18.490 80.750 18.520 ;
        RECT 33.390 18.450 39.800 18.490 ;
        RECT 40.610 18.450 80.750 18.490 ;
        RECT 84.330 17.240 92.560 18.520 ;
      LAYER met3 ;
        RECT 84.280 17.265 92.610 21.995 ;
        RECT 88.150 1.060 89.050 17.265 ;
        RECT 88.110 0.980 90.060 1.060 ;
        RECT 88.110 0.130 90.190 0.980 ;
        RECT 88.150 0.100 89.050 0.130 ;
      LAYER met4 ;
        RECT 44.490 8.685 77.980 39.485 ;
        RECT 84.325 17.285 92.565 21.975 ;
        RECT 88.155 1.000 90.015 1.060 ;
        RECT 88.150 0.100 94.750 1.000 ;
        RECT 93.850 0.000 94.750 0.100 ;
      LAYER met5 ;
        RECT 76.490 21.140 78.090 39.490 ;
        RECT 84.210 21.140 92.680 22.090 ;
        RECT 76.490 17.770 92.680 21.140 ;
        RECT 76.490 8.680 78.090 17.770 ;
        RECT 84.210 17.170 92.680 17.770 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.500000 ;
    PORT
      LAYER li1 ;
        RECT 28.285 32.620 28.615 32.790 ;
        RECT 28.875 32.620 29.205 32.790 ;
        RECT 101.790 21.560 102.290 21.730 ;
        RECT 101.790 18.010 102.290 18.180 ;
        RECT 28.285 17.070 28.615 17.240 ;
        RECT 28.875 17.070 29.205 17.240 ;
      LAYER met1 ;
        RECT 28.150 32.900 30.630 32.910 ;
        RECT 28.150 32.620 30.650 32.900 ;
        RECT 28.305 32.590 28.595 32.620 ;
        RECT 28.895 32.590 29.185 32.620 ;
        RECT 30.280 26.960 30.650 32.620 ;
        RECT 12.700 26.440 13.300 26.560 ;
        RECT 9.550 26.430 13.300 26.440 ;
        RECT 9.550 25.430 13.510 26.430 ;
        RECT 30.140 25.600 30.740 26.960 ;
        RECT 9.550 25.180 13.300 25.430 ;
        RECT 9.550 25.080 13.220 25.180 ;
        RECT 30.280 17.280 30.650 25.600 ;
        RECT 101.520 21.520 102.530 21.980 ;
        RECT 101.810 17.980 102.270 18.210 ;
        RECT 28.220 16.900 30.700 17.280 ;
      LAYER met2 ;
        RECT 9.600 25.030 10.960 26.490 ;
        RECT 12.750 26.430 13.250 26.610 ;
        RECT 30.190 26.430 30.690 27.010 ;
        RECT 12.750 25.750 30.690 26.430 ;
        RECT 12.750 25.130 13.250 25.750 ;
        RECT 30.190 25.550 30.690 25.750 ;
        RECT 101.570 21.470 102.480 22.030 ;
      LAYER met3 ;
        RECT 9.550 25.055 11.010 26.465 ;
        RECT 101.520 21.495 102.530 22.005 ;
        RECT 96.710 4.210 102.550 4.230 ;
        RECT 14.925 4.120 15.815 4.145 ;
        RECT 9.600 3.220 15.930 4.120 ;
        RECT 14.925 3.195 15.815 3.220 ;
        RECT 96.710 3.200 102.560 4.210 ;
        RECT 96.720 3.190 101.530 3.200 ;
      LAYER met4 ;
        RECT 9.595 25.075 10.965 26.445 ;
        RECT 9.630 4.125 10.530 25.075 ;
        RECT 101.565 21.515 102.485 21.985 ;
        RECT 101.570 4.195 102.470 21.515 ;
        RECT 9.625 3.215 10.535 4.125 ;
        RECT 96.765 4.120 97.745 4.145 ;
        RECT 14.920 3.220 97.745 4.120 ;
        RECT 101.535 3.245 102.515 4.195 ;
        RECT 74.530 0.000 75.430 3.220 ;
        RECT 96.765 3.195 97.745 3.220 ;
        RECT 101.570 3.200 102.470 3.245 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.500000 ;
    PORT
      LAYER li1 ;
        RECT 25.435 32.620 25.765 32.790 ;
        RECT 26.025 32.620 26.355 32.790 ;
        RECT 99.335 21.560 99.835 21.730 ;
        RECT 99.335 18.010 99.835 18.180 ;
        RECT 25.435 17.070 25.765 17.240 ;
        RECT 26.025 17.070 26.355 17.240 ;
      LAYER met1 ;
        RECT 23.570 32.900 23.970 32.940 ;
        RECT 23.570 32.580 26.450 32.900 ;
        RECT 11.950 20.850 13.720 22.640 ;
        RECT 23.570 22.200 23.970 32.580 ;
        RECT 23.400 21.010 24.100 22.200 ;
        RECT 99.040 21.520 100.030 21.940 ;
        RECT 11.930 19.270 13.730 20.850 ;
        RECT 11.950 19.230 13.720 19.270 ;
        RECT 23.570 17.280 23.970 21.010 ;
        RECT 99.355 17.980 99.815 18.210 ;
        RECT 23.570 16.980 26.420 17.280 ;
        RECT 23.570 16.930 23.970 16.980 ;
      LAYER met2 ;
        RECT 12.500 22.090 13.100 22.380 ;
        RECT 23.450 22.090 24.050 22.250 ;
        RECT 12.500 21.190 24.050 22.090 ;
        RECT 99.090 21.470 99.980 21.990 ;
        RECT 12.500 21.090 13.100 21.190 ;
        RECT 23.450 20.960 24.050 21.190 ;
        RECT 11.980 19.220 13.680 20.900 ;
      LAYER met3 ;
        RECT 99.040 21.495 100.030 21.965 ;
        RECT 11.930 19.245 13.730 20.875 ;
        RECT 68.980 2.340 72.000 2.430 ;
        RECT 79.510 2.340 82.530 2.430 ;
        RECT 68.980 1.440 82.530 2.340 ;
        RECT 68.980 1.400 72.000 1.440 ;
        RECT 79.510 1.400 82.530 1.440 ;
      LAYER met4 ;
        RECT 99.080 21.945 99.980 22.090 ;
        RECT 99.080 21.515 99.985 21.945 ;
        RECT 11.975 19.265 13.685 20.855 ;
        RECT 12.290 2.340 13.190 19.265 ;
        RECT 69.025 2.340 71.955 2.435 ;
        RECT 12.290 1.440 71.955 2.340 ;
        RECT 55.210 0.000 56.110 1.440 ;
        RECT 69.025 1.395 71.955 1.440 ;
        RECT 79.555 2.340 82.485 2.435 ;
        RECT 99.080 2.340 99.980 21.515 ;
        RECT 79.555 1.440 99.980 2.340 ;
        RECT 79.555 1.395 82.485 1.440 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 101.610 80.140 108.570 84.330 ;
        RECT 122.870 76.790 126.940 80.980 ;
        RECT 113.950 64.950 116.060 70.140 ;
        RECT 120.250 69.090 147.210 72.280 ;
        RECT 124.410 66.085 126.590 67.690 ;
        RECT 128.620 66.125 131.760 67.730 ;
        RECT 111.750 60.490 114.710 63.680 ;
        RECT 94.970 56.850 95.810 56.870 ;
        RECT 94.970 55.265 97.520 56.850 ;
        RECT 95.760 55.245 97.520 55.265 ;
        RECT 124.570 53.890 139.140 64.080 ;
        RECT 31.810 21.460 43.500 38.650 ;
        RECT 100.800 26.765 103.260 26.780 ;
        RECT 98.385 22.590 103.260 26.765 ;
        RECT 98.385 22.575 100.845 22.590 ;
        RECT 39.870 17.460 43.500 21.460 ;
        RECT 104.860 19.940 110.480 26.780 ;
      LAYER li1 ;
        RECT 101.790 83.980 108.390 84.150 ;
        RECT 98.900 80.890 100.310 83.050 ;
        RECT 101.790 80.490 101.960 83.980 ;
        RECT 107.650 82.190 107.820 83.255 ;
        RECT 108.220 82.190 108.390 83.980 ;
        RECT 107.650 81.880 108.400 82.190 ;
        RECT 107.650 81.215 107.820 81.880 ;
        RECT 108.220 80.490 108.390 81.880 ;
        RECT 101.790 80.320 108.390 80.490 ;
        RECT 123.050 80.630 126.760 80.800 ;
        RECT 123.050 77.140 123.220 80.630 ;
        RECT 124.100 77.865 124.270 79.905 ;
        RECT 125.060 77.865 125.230 79.905 ;
        RECT 126.020 77.865 126.190 79.905 ;
        RECT 126.590 79.870 126.760 80.630 ;
        RECT 126.590 79.140 126.840 79.870 ;
        RECT 126.590 77.140 126.760 79.140 ;
        RECT 132.865 78.545 134.275 80.705 ;
        RECT 123.050 76.970 126.760 77.140 ;
        RECT 120.430 71.930 147.030 72.100 ;
        RECT 114.130 69.790 115.880 69.960 ;
        RECT 114.130 65.300 114.300 69.790 ;
        RECT 115.140 67.050 115.310 69.065 ;
        RECT 115.710 67.050 115.880 69.790 ;
        RECT 120.430 69.440 120.600 71.930 ;
        RECT 146.290 70.760 146.460 71.205 ;
        RECT 146.860 70.760 147.030 71.930 ;
        RECT 146.290 70.380 147.030 70.760 ;
        RECT 146.290 70.165 146.460 70.380 ;
        RECT 146.860 69.440 147.030 70.380 ;
        RECT 120.430 69.270 147.030 69.440 ;
        RECT 124.600 67.415 126.400 67.585 ;
        RECT 128.810 67.455 131.570 67.625 ;
        RECT 115.120 66.180 115.920 67.050 ;
        RECT 124.940 66.275 125.150 67.415 ;
        RECT 126.025 66.250 126.315 67.415 ;
        RECT 128.895 66.290 129.185 67.455 ;
        RECT 129.430 66.995 129.700 67.455 ;
        RECT 130.380 66.655 130.890 67.455 ;
        RECT 115.140 66.025 115.310 66.180 ;
        RECT 115.710 65.300 115.880 66.180 ;
        RECT 114.130 65.130 115.880 65.300 ;
        RECT 126.530 63.900 127.230 63.930 ;
        RECT 124.750 63.730 138.960 63.900 ;
        RECT 111.930 63.330 114.530 63.500 ;
        RECT 111.930 60.840 112.100 63.330 ;
        RECT 113.790 62.430 113.960 62.605 ;
        RECT 114.360 62.430 114.530 63.330 ;
        RECT 113.770 62.060 114.530 62.430 ;
        RECT 113.790 61.565 113.960 62.060 ;
        RECT 114.360 60.840 114.530 62.060 ;
        RECT 111.930 60.670 114.530 60.840 ;
        RECT 95.160 56.595 95.620 56.765 ;
        RECT 95.245 55.430 95.535 56.595 ;
        RECT 95.950 56.575 97.330 56.745 ;
        RECT 96.290 55.435 96.500 56.575 ;
        RECT 124.750 54.240 124.920 63.730 ;
        RECT 126.610 54.965 126.780 63.005 ;
        RECT 129.190 54.965 129.360 63.005 ;
        RECT 131.770 54.965 131.940 63.005 ;
        RECT 134.350 54.965 134.520 63.005 ;
        RECT 136.930 54.965 137.100 63.005 ;
        RECT 138.790 54.240 138.960 63.730 ;
        RECT 124.750 54.070 138.960 54.240 ;
        RECT 33.380 38.470 34.320 38.710 ;
        RECT 37.250 38.470 38.190 38.670 ;
        RECT 41.080 38.470 42.020 38.700 ;
        RECT 31.990 38.300 35.660 38.470 ;
        RECT 14.890 33.890 15.240 36.050 ;
        RECT 31.990 21.810 32.160 38.300 ;
        RECT 33.380 38.290 34.320 38.300 ;
        RECT 32.560 22.535 32.730 37.575 ;
        RECT 33.740 22.535 33.910 37.575 ;
        RECT 34.920 22.535 35.090 37.575 ;
        RECT 35.490 21.810 35.660 38.300 ;
        RECT 31.990 21.640 35.660 21.810 ;
        RECT 36.020 38.300 39.690 38.470 ;
        RECT 36.020 21.810 36.190 38.300 ;
        RECT 37.250 38.250 38.190 38.300 ;
        RECT 36.590 22.535 36.760 37.575 ;
        RECT 37.770 22.535 37.940 37.575 ;
        RECT 38.950 22.535 39.120 37.575 ;
        RECT 39.520 21.810 39.690 38.300 ;
        RECT 36.020 21.640 39.690 21.810 ;
        RECT 40.050 38.300 43.320 38.470 ;
        RECT 40.050 17.810 40.220 38.300 ;
        RECT 41.080 38.280 42.020 38.300 ;
        RECT 40.620 18.535 40.790 37.575 ;
        RECT 41.600 18.535 41.770 37.575 ;
        RECT 42.580 18.535 42.750 37.575 ;
        RECT 43.150 17.810 43.320 38.300 ;
        RECT 96.120 28.290 96.810 30.450 ;
        RECT 97.900 27.240 115.800 28.590 ;
        RECT 99.350 26.585 99.850 27.240 ;
        RECT 100.450 26.600 101.150 26.640 ;
        RECT 101.800 26.600 102.300 27.240 ;
        RECT 107.600 26.600 108.100 27.240 ;
        RECT 100.450 26.590 103.080 26.600 ;
        RECT 100.400 26.585 103.080 26.590 ;
        RECT 98.565 26.440 103.080 26.585 ;
        RECT 98.565 26.415 100.665 26.440 ;
        RECT 98.565 25.690 98.735 26.415 ;
        RECT 98.550 25.340 99.350 25.690 ;
        RECT 98.565 22.925 98.735 25.340 ;
        RECT 99.135 23.650 99.305 25.340 ;
        RECT 100.495 22.925 100.665 26.415 ;
        RECT 98.565 22.755 100.665 22.925 ;
        RECT 100.980 26.430 103.080 26.440 ;
        RECT 100.980 22.940 101.150 26.430 ;
        RECT 102.340 25.690 102.510 25.705 ;
        RECT 102.910 25.690 103.080 26.430 ;
        RECT 105.040 26.430 110.300 26.600 ;
        RECT 105.040 25.690 105.210 26.430 ;
        RECT 105.580 25.710 105.810 26.430 ;
        RECT 107.160 25.710 107.390 26.430 ;
        RECT 108.740 25.710 108.970 26.430 ;
        RECT 102.290 25.240 105.210 25.690 ;
        RECT 102.340 23.665 102.510 25.240 ;
        RECT 102.910 22.940 103.080 25.240 ;
        RECT 100.980 22.770 103.080 22.940 ;
        RECT 105.040 20.290 105.210 25.240 ;
        RECT 105.610 21.020 105.780 25.710 ;
        RECT 107.190 21.020 107.360 25.710 ;
        RECT 108.770 21.020 108.940 25.710 ;
        RECT 110.130 20.290 110.300 26.430 ;
        RECT 105.040 20.120 110.300 20.290 ;
        RECT 40.050 17.640 43.320 17.810 ;
      LAYER met1 ;
        RECT 108.670 84.950 109.850 86.020 ;
        RECT 107.620 83.230 107.850 83.235 ;
        RECT 98.960 83.020 100.350 83.070 ;
        RECT 98.950 81.000 100.350 83.020 ;
        RECT 107.560 81.260 107.930 83.230 ;
        RECT 108.120 81.940 108.520 82.650 ;
        RECT 107.620 81.235 107.850 81.260 ;
        RECT 98.950 80.915 100.260 81.000 ;
        RECT 132.915 80.670 134.225 80.675 ;
        RECT 124.070 78.520 124.300 79.885 ;
        RECT 124.000 78.000 124.370 78.520 ;
        RECT 125.030 78.510 125.260 79.885 ;
        RECT 125.990 78.530 126.220 79.885 ;
        RECT 126.560 79.640 126.870 79.930 ;
        RECT 126.540 79.140 126.980 79.640 ;
        RECT 126.560 79.080 126.870 79.140 ;
        RECT 132.890 78.560 134.230 80.670 ;
        RECT 124.070 77.885 124.300 78.000 ;
        RECT 124.950 77.990 125.320 78.510 ;
        RECT 125.910 78.010 126.280 78.530 ;
        RECT 125.030 77.885 125.260 77.990 ;
        RECT 125.990 77.885 126.220 78.010 ;
        RECT 146.260 71.160 146.490 71.185 ;
        RECT 146.190 70.230 146.550 71.160 ;
        RECT 146.260 70.185 146.490 70.230 ;
        RECT 115.110 67.010 115.340 69.045 ;
        RECT 129.120 67.780 129.710 67.970 ;
        RECT 124.600 67.720 126.400 67.740 ;
        RECT 124.560 67.270 126.400 67.720 ;
        RECT 128.810 67.300 131.570 67.780 ;
        RECT 124.600 67.260 126.400 67.270 ;
        RECT 115.050 66.220 115.620 67.010 ;
        RECT 115.110 66.045 115.340 66.220 ;
        RECT 126.480 63.960 127.270 64.080 ;
        RECT 126.470 63.710 127.290 63.960 ;
        RECT 113.760 62.510 113.990 62.585 ;
        RECT 113.730 62.170 114.160 62.510 ;
        RECT 113.760 61.585 113.990 62.170 ;
        RECT 126.580 61.940 126.810 62.985 ;
        RECT 129.160 61.940 129.390 62.985 ;
        RECT 131.740 62.010 131.970 62.985 ;
        RECT 126.580 60.720 126.850 61.940 ;
        RECT 129.160 60.720 129.430 61.940 ;
        RECT 131.740 60.790 132.000 62.010 ;
        RECT 134.320 61.900 134.550 62.985 ;
        RECT 126.580 57.280 126.810 60.720 ;
        RECT 95.160 56.840 95.620 56.920 ;
        RECT 95.920 56.900 96.390 56.960 ;
        RECT 126.470 56.950 126.850 57.280 ;
        RECT 129.160 57.050 129.390 60.720 ;
        RECT 95.920 56.840 97.330 56.900 ;
        RECT 94.880 56.420 97.330 56.840 ;
        RECT 126.460 55.960 126.940 56.950 ;
        RECT 128.990 56.000 129.610 57.050 ;
        RECT 131.740 56.980 131.970 60.790 ;
        RECT 134.320 60.680 134.580 61.900 ;
        RECT 134.320 57.030 134.550 60.680 ;
        RECT 136.900 57.050 137.130 62.985 ;
        RECT 126.580 54.985 126.810 55.960 ;
        RECT 129.160 54.985 129.390 56.000 ;
        RECT 131.610 55.930 132.230 56.980 ;
        RECT 134.130 55.980 134.750 57.030 ;
        RECT 136.720 56.000 137.340 57.050 ;
        RECT 131.740 54.985 131.970 55.930 ;
        RECT 134.320 54.985 134.550 55.980 ;
        RECT 136.900 54.985 137.130 56.000 ;
        RECT 0.970 43.960 2.980 48.190 ;
        RECT 0.970 43.290 104.820 43.960 ;
        RECT 0.960 42.380 104.820 43.290 ;
        RECT 0.960 42.270 2.980 42.380 ;
        RECT 0.960 40.550 2.970 42.270 ;
        RECT 0.960 38.730 42.020 40.550 ;
        RECT 0.960 38.250 42.080 38.730 ;
        RECT 0.960 38.230 42.020 38.250 ;
        RECT 0.960 37.370 2.970 38.230 ;
        RECT 14.640 35.790 15.530 38.230 ;
        RECT 37.190 38.220 38.250 38.230 ;
        RECT 32.530 36.500 32.760 37.555 ;
        RECT 33.710 36.510 33.940 37.555 ;
        RECT 14.830 35.700 15.310 35.790 ;
        RECT 32.350 35.770 32.890 36.500 ;
        RECT 33.560 35.780 34.100 36.510 ;
        RECT 34.890 36.480 35.120 37.555 ;
        RECT 14.940 33.915 15.190 35.700 ;
        RECT 32.530 22.555 32.760 35.770 ;
        RECT 33.710 22.555 33.940 35.780 ;
        RECT 34.740 35.750 35.280 36.480 ;
        RECT 36.560 36.460 36.790 37.555 ;
        RECT 34.890 22.555 35.120 35.750 ;
        RECT 36.380 35.730 36.920 36.460 ;
        RECT 37.740 36.410 37.970 37.555 ;
        RECT 36.560 22.555 36.790 35.730 ;
        RECT 37.580 35.680 38.120 36.410 ;
        RECT 38.920 36.380 39.150 37.555 ;
        RECT 40.590 36.380 40.820 37.555 ;
        RECT 41.570 36.400 41.800 37.555 ;
        RECT 42.550 36.420 42.780 37.555 ;
        RECT 37.740 22.555 37.970 35.680 ;
        RECT 38.770 35.650 39.310 36.380 ;
        RECT 40.380 35.650 40.920 36.380 ;
        RECT 41.450 35.690 41.920 36.400 ;
        RECT 42.430 35.710 42.900 36.420 ;
        RECT 38.920 22.555 39.150 35.650 ;
        RECT 40.590 18.555 40.820 35.650 ;
        RECT 41.570 18.555 41.800 35.690 ;
        RECT 42.550 18.555 42.780 35.710 ;
        RECT 96.170 28.590 96.760 30.420 ;
        RECT 96.100 28.270 99.950 28.590 ;
        RECT 97.750 28.260 99.950 28.270 ;
        RECT 103.240 27.240 104.820 42.380 ;
        RECT 99.105 23.670 99.335 25.670 ;
        RECT 102.310 23.685 102.540 25.685 ;
        RECT 105.580 21.040 105.810 26.040 ;
        RECT 107.160 21.040 107.390 26.040 ;
        RECT 108.740 21.040 108.970 26.040 ;
      LAYER met2 ;
        RECT 108.720 85.930 109.800 86.070 ;
        RECT 108.720 84.890 109.850 85.930 ;
        RECT 99.010 80.950 100.300 83.120 ;
        RECT 107.610 82.840 107.880 83.280 ;
        RECT 107.600 81.920 107.950 82.840 ;
        RECT 108.220 82.700 108.570 82.800 ;
        RECT 107.610 81.210 107.880 81.920 ;
        RECT 108.170 81.890 108.570 82.700 ;
        RECT 108.220 81.880 108.570 81.890 ;
        RECT 126.590 79.090 126.930 79.690 ;
        RECT 124.000 78.600 124.370 78.640 ;
        RECT 124.000 77.940 126.330 78.600 ;
        RECT 132.920 78.560 134.180 80.730 ;
        RECT 132.940 78.510 134.180 78.560 ;
        RECT 124.000 77.910 124.370 77.940 ;
        RECT 146.240 70.960 146.500 71.210 ;
        RECT 146.240 70.400 146.570 70.960 ;
        RECT 146.240 70.180 146.500 70.400 ;
        RECT 129.190 68.020 129.760 68.050 ;
        RECT 124.610 67.220 125.030 67.770 ;
        RECT 129.170 67.500 129.760 68.020 ;
        RECT 129.190 67.480 129.760 67.500 ;
        RECT 115.120 67.060 115.570 67.080 ;
        RECT 115.100 66.170 115.570 67.060 ;
        RECT 115.120 66.130 115.570 66.170 ;
        RECT 126.530 63.690 127.220 64.130 ;
        RECT 113.780 62.120 114.170 62.560 ;
        RECT 126.470 57.010 126.850 57.280 ;
        RECT 129.040 57.010 129.560 57.100 ;
        RECT 131.660 57.010 132.180 57.030 ;
        RECT 134.180 57.010 134.700 57.080 ;
        RECT 136.770 57.020 137.290 57.100 ;
        RECT 136.260 57.010 137.810 57.020 ;
        RECT 95.530 56.960 96.390 56.970 ;
        RECT 95.520 56.210 96.440 56.960 ;
        RECT 126.160 56.950 137.830 57.010 ;
        RECT 95.530 56.180 96.390 56.210 ;
        RECT 126.040 55.990 137.830 56.950 ;
        RECT 126.160 55.940 137.830 55.990 ;
        RECT 126.510 55.910 126.890 55.940 ;
        RECT 131.660 55.880 132.180 55.940 ;
        RECT 134.180 55.930 134.700 55.940 ;
        RECT 136.260 55.730 137.810 55.940 ;
        RECT 1.020 43.340 2.930 48.240 ;
        RECT 1.010 42.220 2.930 43.340 ;
        RECT 1.010 37.320 2.920 42.220 ;
        RECT 33.380 38.240 34.320 38.760 ;
        RECT 32.400 36.350 32.840 36.550 ;
        RECT 33.540 36.350 34.170 38.240 ;
        RECT 37.250 38.200 38.190 38.720 ;
        RECT 41.080 38.230 42.020 38.750 ;
        RECT 34.790 36.350 35.230 36.530 ;
        RECT 36.430 36.350 36.870 36.510 ;
        RECT 37.430 36.460 38.060 38.200 ;
        RECT 37.430 36.350 38.070 36.460 ;
        RECT 38.820 36.350 39.260 36.430 ;
        RECT 40.430 36.350 40.870 36.430 ;
        RECT 41.260 36.350 41.890 38.230 ;
        RECT 42.480 36.350 42.850 36.470 ;
        RECT 32.400 35.750 42.850 36.350 ;
        RECT 32.400 35.720 32.840 35.750 ;
        RECT 33.610 35.730 34.050 35.750 ;
        RECT 34.790 35.700 35.230 35.750 ;
        RECT 36.430 35.680 36.870 35.750 ;
        RECT 37.630 35.630 38.070 35.750 ;
        RECT 38.820 35.600 39.260 35.750 ;
        RECT 40.430 35.600 40.870 35.750 ;
        RECT 41.500 35.640 41.870 35.750 ;
        RECT 42.480 35.660 42.850 35.750 ;
      LAYER met3 ;
        RECT 1.020 86.290 2.940 88.780 ;
        RECT 9.870 86.290 14.140 86.300 ;
        RECT 1.020 84.860 14.140 86.290 ;
        RECT 108.670 84.925 109.850 86.045 ;
        RECT 1.020 82.410 2.940 84.860 ;
        RECT 99.050 81.035 100.340 82.965 ;
        RECT 107.550 82.810 108.000 82.815 ;
        RECT 107.550 82.775 108.560 82.810 ;
        RECT 107.550 81.945 108.620 82.775 ;
        RECT 107.600 81.905 108.620 81.945 ;
        RECT 107.600 81.870 108.560 81.905 ;
        RECT 126.540 79.115 126.980 79.665 ;
        RECT 123.950 77.935 124.420 78.615 ;
        RECT 132.870 78.585 134.230 80.705 ;
        RECT 146.220 70.450 146.710 70.940 ;
        RECT 146.220 70.425 146.620 70.450 ;
        RECT 124.560 67.245 125.080 67.745 ;
        RECT 129.140 67.505 129.810 68.025 ;
        RECT 115.070 66.155 115.620 67.055 ;
        RECT 113.770 62.060 114.380 65.570 ;
        RECT 126.480 63.715 127.270 64.105 ;
        RECT 126.470 56.975 126.850 57.280 ;
        RECT 95.480 56.205 96.440 56.945 ;
        RECT 126.460 55.935 126.940 56.975 ;
        RECT 0.970 43.315 2.980 48.215 ;
        RECT 0.960 42.245 2.980 43.315 ;
        RECT 0.960 37.345 2.970 42.245 ;
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
        RECT 11.295 86.080 14.005 86.145 ;
        RECT 98.900 86.090 100.390 86.110 ;
        RECT 98.550 86.080 109.690 86.090 ;
        RECT 11.290 86.025 109.690 86.080 ;
        RECT 11.290 85.800 109.805 86.025 ;
        RECT 110.230 85.800 111.390 85.850 ;
        RECT 122.570 85.800 124.370 85.840 ;
        RECT 11.290 85.350 124.370 85.800 ;
        RECT 11.290 85.050 124.390 85.350 ;
        RECT 11.290 85.040 123.080 85.050 ;
        RECT 11.290 85.030 113.710 85.040 ;
        RECT 114.350 85.030 123.080 85.040 ;
        RECT 11.290 85.010 109.805 85.030 ;
        RECT 11.290 84.940 100.390 85.010 ;
        RECT 108.715 84.945 109.805 85.010 ;
        RECT 11.295 84.915 14.005 84.940 ;
        RECT 95.520 56.925 96.290 84.940 ;
        RECT 98.900 80.890 100.390 84.940 ;
        RECT 110.230 82.810 111.390 85.030 ;
        RECT 124.040 82.810 124.390 85.050 ;
        RECT 129.190 82.810 129.780 82.920 ;
        RECT 133.870 82.810 135.860 82.820 ;
        RECT 146.250 82.810 146.740 82.880 ;
        RECT 107.580 81.960 111.450 82.810 ;
        RECT 123.640 82.220 146.740 82.810 ;
        RECT 107.590 81.950 108.770 81.960 ;
        RECT 107.590 81.925 108.575 81.950 ;
        RECT 107.590 81.910 108.570 81.925 ;
        RECT 110.230 65.580 111.390 81.960 ;
        RECT 124.080 78.595 124.470 82.220 ;
        RECT 126.490 81.980 127.210 82.220 ;
        RECT 123.995 77.955 124.470 78.595 ;
        RECT 124.080 68.360 124.470 77.955 ;
        RECT 124.060 67.750 124.470 68.360 ;
        RECT 124.060 67.740 125.010 67.750 ;
        RECT 124.060 67.320 125.070 67.740 ;
        RECT 124.440 67.280 125.070 67.320 ;
        RECT 124.605 67.265 125.035 67.280 ;
        RECT 115.090 67.035 115.390 67.120 ;
        RECT 115.090 66.175 115.575 67.035 ;
        RECT 115.090 65.580 115.390 66.175 ;
        RECT 110.230 64.820 115.820 65.580 ;
        RECT 126.510 65.510 127.200 81.980 ;
        RECT 129.190 68.005 129.780 82.220 ;
        RECT 132.840 82.190 135.860 82.220 ;
        RECT 132.840 78.630 134.220 82.190 ;
        RECT 132.915 78.605 134.185 78.630 ;
        RECT 146.250 70.360 146.740 82.220 ;
        RECT 129.185 67.580 129.780 68.005 ;
        RECT 129.185 67.525 129.765 67.580 ;
        RECT 110.230 64.790 111.390 64.820 ;
        RECT 113.460 64.750 114.380 64.820 ;
        RECT 113.770 62.060 114.380 64.750 ;
        RECT 126.510 64.620 127.220 65.510 ;
        RECT 126.520 64.085 127.220 64.620 ;
        RECT 126.520 63.735 127.225 64.085 ;
        RECT 126.520 57.280 127.220 63.735 ;
        RECT 126.470 56.950 127.220 57.280 ;
        RECT 95.520 56.350 96.395 56.925 ;
        RECT 95.525 56.225 96.395 56.350 ;
        RECT 126.505 55.970 127.220 56.950 ;
        RECT 126.505 55.960 127.200 55.970 ;
        RECT 126.505 55.955 126.895 55.960 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 98.120 83.400 101.090 83.830 ;
        RECT 98.120 77.320 98.550 83.400 ;
        RECT 100.660 77.320 101.090 83.400 ;
        RECT 98.120 76.890 101.090 77.320 ;
        RECT 114.290 71.290 119.290 73.450 ;
        RECT 97.120 67.490 100.090 67.920 ;
        RECT 97.120 61.410 97.550 67.490 ;
        RECT 99.660 61.410 100.090 67.490 ;
        RECT 116.230 65.300 120.200 69.300 ;
        RECT 97.120 60.980 100.090 61.410 ;
        RECT 115.100 59.280 118.590 64.280 ;
        RECT 119.720 59.670 122.580 62.670 ;
        RECT 95.175 54.150 95.605 54.935 ;
        RECT 103.890 53.700 105.900 56.700 ;
        RECT 14.110 36.400 16.020 36.830 ;
        RECT 14.110 12.540 14.540 36.400 ;
        RECT 15.590 12.540 16.020 36.400 ;
        RECT 14.110 12.110 16.020 12.540 ;
        RECT 16.110 36.400 18.020 36.830 ;
        RECT 16.110 12.540 16.540 36.400 ;
        RECT 17.590 12.540 18.020 36.400 ;
        RECT 16.110 12.110 18.020 12.540 ;
        RECT 18.120 36.400 20.030 36.830 ;
        RECT 18.120 12.540 18.550 36.400 ;
        RECT 19.600 12.540 20.030 36.400 ;
        RECT 18.120 12.110 20.030 12.540 ;
        RECT 20.120 36.400 22.030 36.830 ;
        RECT 20.120 12.540 20.550 36.400 ;
        RECT 21.600 12.540 22.030 36.400 ;
        RECT 20.120 12.110 22.030 12.540 ;
        RECT 22.130 36.400 24.040 36.830 ;
        RECT 22.130 12.540 22.560 36.400 ;
        RECT 23.610 12.540 24.040 36.400 ;
        RECT 24.520 16.430 27.270 33.430 ;
        RECT 27.370 16.430 30.120 33.430 ;
        RECT 95.340 30.800 97.590 31.230 ;
        RECT 22.130 12.110 24.040 12.540 ;
        RECT 20.050 9.020 24.200 12.020 ;
        RECT 24.380 8.950 31.110 15.950 ;
        RECT 31.690 8.900 38.420 20.900 ;
        RECT 39.070 16.090 41.320 16.520 ;
        RECT 39.070 9.330 39.500 16.090 ;
        RECT 40.890 9.330 41.320 16.090 ;
        RECT 39.070 8.900 41.320 9.330 ;
        RECT 95.340 7.240 95.770 30.800 ;
        RECT 97.160 7.240 97.590 30.800 ;
        RECT 98.405 17.370 100.765 22.370 ;
        RECT 100.860 17.370 103.220 22.370 ;
        RECT 104.450 19.200 117.310 19.630 ;
        RECT 104.450 18.170 104.880 19.200 ;
        RECT 116.880 18.170 117.310 19.200 ;
        RECT 104.450 17.740 117.310 18.170 ;
        RECT 98.450 9.090 100.810 16.780 ;
        RECT 100.900 9.090 103.260 16.780 ;
        RECT 103.950 11.540 110.260 17.140 ;
        RECT 95.340 6.810 97.590 7.240 ;
      LAYER li1 ;
        RECT 98.250 83.530 100.960 83.700 ;
        RECT 98.250 79.820 98.420 83.530 ;
        RECT 95.500 79.080 98.470 79.820 ;
        RECT 95.520 59.550 96.300 79.080 ;
        RECT 98.250 77.190 98.420 79.080 ;
        RECT 100.790 77.190 100.960 83.530 ;
        RECT 98.250 77.020 100.960 77.190 ;
        RECT 114.420 73.150 119.160 73.320 ;
        RECT 114.420 72.770 114.590 73.150 ;
        RECT 114.200 72.230 114.590 72.770 ;
        RECT 115.380 72.750 118.300 73.150 ;
        RECT 115.270 72.580 118.310 72.750 ;
        RECT 114.420 71.590 114.590 72.230 ;
        RECT 118.990 71.590 119.160 73.150 ;
        RECT 114.420 71.420 119.160 71.590 ;
        RECT 116.360 69.000 120.070 69.170 ;
        RECT 97.250 67.620 99.960 67.790 ;
        RECT 97.250 61.280 97.420 67.620 ;
        RECT 97.790 61.280 98.360 61.350 ;
        RECT 99.790 61.280 99.960 67.620 ;
        RECT 116.360 65.600 116.530 69.000 ;
        RECT 117.410 66.280 117.580 68.320 ;
        RECT 118.370 66.280 118.540 68.320 ;
        RECT 119.330 66.280 119.500 68.320 ;
        RECT 119.900 65.600 120.070 69.000 ;
        RECT 116.360 65.430 120.070 65.600 ;
        RECT 117.310 64.150 117.980 65.430 ;
        RECT 97.250 61.110 99.960 61.280 ;
        RECT 115.230 63.980 118.460 64.150 ;
        RECT 97.790 59.550 98.360 61.110 ;
        RECT 95.520 59.010 98.360 59.550 ;
        RECT 115.230 59.580 115.400 63.980 ;
        RECT 116.280 60.260 116.450 63.300 ;
        RECT 117.240 60.260 117.410 63.300 ;
        RECT 118.290 60.760 118.460 63.980 ;
        RECT 119.850 62.370 122.450 62.540 ;
        RECT 119.850 60.760 120.020 62.370 ;
        RECT 118.290 60.210 120.070 60.760 ;
        RECT 121.710 60.650 121.880 61.690 ;
        RECT 118.290 59.580 118.460 60.210 ;
        RECT 119.850 59.970 120.020 60.210 ;
        RECT 122.280 59.970 122.450 62.370 ;
        RECT 119.850 59.800 122.450 59.970 ;
        RECT 119.950 59.640 120.840 59.800 ;
        RECT 115.230 59.410 118.460 59.580 ;
        RECT 95.550 58.970 98.360 59.010 ;
        RECT 95.245 54.045 95.535 54.770 ;
        RECT 95.160 53.875 95.620 54.045 ;
        RECT 96.270 54.025 96.500 54.845 ;
        RECT 97.790 54.720 98.360 58.970 ;
        RECT 104.020 56.400 105.770 56.570 ;
        RECT 104.020 54.720 104.190 56.400 ;
        RECT 97.790 54.190 104.200 54.720 ;
        RECT 105.030 54.680 105.200 55.720 ;
        RECT 97.790 54.030 98.360 54.190 ;
        RECT 97.100 54.025 98.360 54.030 ;
        RECT 95.950 53.855 98.360 54.025 ;
        RECT 97.100 53.850 98.360 53.855 ;
        RECT 104.020 54.000 104.190 54.190 ;
        RECT 105.600 54.000 105.770 56.400 ;
        RECT 104.020 53.830 105.770 54.000 ;
        RECT 14.240 36.530 15.890 36.700 ;
        RECT 14.240 12.410 14.410 36.530 ;
        RECT 15.720 12.410 15.890 36.530 ;
        RECT 16.240 36.530 17.890 36.700 ;
        RECT 16.240 12.410 16.410 36.530 ;
        RECT 17.720 12.410 17.890 36.530 ;
        RECT 18.250 36.530 19.900 36.700 ;
        RECT 18.250 12.410 18.420 36.530 ;
        RECT 19.730 12.410 19.900 36.530 ;
        RECT 20.250 36.530 21.900 36.700 ;
        RECT 20.250 12.410 20.420 36.530 ;
        RECT 21.730 12.410 21.900 36.530 ;
        RECT 22.260 36.530 23.910 36.700 ;
        RECT 22.260 12.410 22.430 36.530 ;
        RECT 23.740 12.410 23.910 36.530 ;
        RECT 24.650 33.130 27.140 33.300 ;
        RECT 24.650 16.730 24.820 33.130 ;
        RECT 26.970 16.750 27.140 33.130 ;
        RECT 27.500 33.130 29.990 33.300 ;
        RECT 27.500 16.750 27.670 33.130 ;
        RECT 26.300 16.730 28.050 16.750 ;
        RECT 29.820 16.730 29.990 33.130 ;
        RECT 95.470 30.930 97.460 31.100 ;
        RECT 24.650 16.560 29.990 16.730 ;
        RECT 31.820 20.600 38.290 20.770 ;
        RECT 26.300 16.190 28.050 16.560 ;
        RECT 14.240 12.240 23.910 12.410 ;
        RECT 24.510 15.650 30.980 15.820 ;
        RECT 15.080 11.890 22.770 12.240 ;
        RECT 15.080 11.720 24.070 11.890 ;
        RECT 20.180 9.320 20.350 11.720 ;
        RECT 20.750 10.000 20.920 11.040 ;
        RECT 23.330 10.000 23.500 11.040 ;
        RECT 21.310 9.320 22.960 9.400 ;
        RECT 23.900 9.320 24.070 11.720 ;
        RECT 20.180 9.150 24.070 9.320 ;
        RECT 24.510 9.250 24.680 15.650 ;
        RECT 25.080 9.930 25.250 14.970 ;
        RECT 27.660 9.930 27.830 14.970 ;
        RECT 30.240 9.930 30.410 14.970 ;
        RECT 26.880 9.250 28.070 9.270 ;
        RECT 30.810 9.250 30.980 15.650 ;
        RECT 21.310 8.960 22.960 9.150 ;
        RECT 24.510 9.080 30.980 9.250 ;
        RECT 31.820 9.200 31.990 20.600 ;
        RECT 32.390 9.880 32.560 19.920 ;
        RECT 34.970 9.880 35.140 19.920 ;
        RECT 37.550 9.880 37.720 19.920 ;
        RECT 34.080 9.200 35.500 9.240 ;
        RECT 38.120 9.200 38.290 20.600 ;
        RECT 26.880 8.780 28.070 9.080 ;
        RECT 31.820 9.030 38.290 9.200 ;
        RECT 39.200 16.220 41.190 16.390 ;
        RECT 39.200 9.200 39.370 16.220 ;
        RECT 41.020 9.200 41.190 16.220 ;
        RECT 39.200 9.030 41.190 9.200 ;
        RECT 34.080 8.830 35.500 9.030 ;
        RECT 39.600 8.540 40.480 9.030 ;
        RECT 95.470 7.110 95.640 30.930 ;
        RECT 97.290 8.110 97.460 30.930 ;
        RECT 100.395 22.240 101.220 22.245 ;
        RECT 98.535 22.070 103.090 22.240 ;
        RECT 98.535 17.670 98.705 22.070 ;
        RECT 100.465 17.670 100.635 22.070 ;
        RECT 100.990 17.670 101.160 22.070 ;
        RECT 102.920 17.670 103.090 22.070 ;
        RECT 104.580 19.330 117.180 19.500 ;
        RECT 104.580 18.040 104.750 19.330 ;
        RECT 117.010 18.040 117.180 19.330 ;
        RECT 104.580 17.870 117.180 18.040 ;
        RECT 98.535 17.500 103.090 17.670 ;
        RECT 100.150 17.495 101.215 17.500 ;
        RECT 100.150 16.650 100.550 17.495 ;
        RECT 100.750 17.440 100.960 17.495 ;
        RECT 105.250 17.010 105.550 17.870 ;
        RECT 104.080 16.840 110.130 17.010 ;
        RECT 98.580 16.480 100.680 16.650 ;
        RECT 98.580 10.890 98.750 16.480 ;
        RECT 99.150 10.890 99.320 16.110 ;
        RECT 98.580 10.390 99.320 10.890 ;
        RECT 98.580 9.390 98.750 10.390 ;
        RECT 99.150 10.070 99.320 10.390 ;
        RECT 100.510 9.390 100.680 16.480 ;
        RECT 101.030 16.480 103.130 16.650 ;
        RECT 101.030 9.390 101.200 16.480 ;
        RECT 102.390 10.940 102.560 16.110 ;
        RECT 102.960 10.940 103.130 16.480 ;
        RECT 104.080 13.940 104.250 16.840 ;
        RECT 103.650 13.690 104.250 13.940 ;
        RECT 102.390 10.790 103.200 10.940 ;
        RECT 103.650 10.790 103.850 13.690 ;
        RECT 104.080 11.840 104.250 13.690 ;
        RECT 104.650 11.840 104.820 16.160 ;
        RECT 106.230 11.840 106.400 16.160 ;
        RECT 107.810 11.840 107.980 16.160 ;
        RECT 109.390 11.840 109.560 16.160 ;
        RECT 109.960 11.840 110.130 16.840 ;
        RECT 104.080 11.670 110.130 11.840 ;
        RECT 102.390 10.590 103.850 10.790 ;
        RECT 102.390 10.440 103.200 10.590 ;
        RECT 102.390 10.070 102.560 10.440 ;
        RECT 102.960 9.390 103.130 10.440 ;
        RECT 98.580 9.220 103.130 9.390 ;
        RECT 100.300 9.190 101.450 9.220 ;
        RECT 100.400 8.890 101.350 9.190 ;
        RECT 106.600 8.890 107.400 11.670 ;
        RECT 97.290 8.100 97.830 8.110 ;
        RECT 98.400 8.100 111.900 8.890 ;
        RECT 97.290 7.740 111.900 8.100 ;
        RECT 97.290 7.110 97.460 7.740 ;
        RECT 98.400 7.290 111.900 7.740 ;
        RECT 95.470 6.940 97.460 7.110 ;
      LAYER met1 ;
        RECT 114.170 72.770 114.580 72.830 ;
        RECT 114.150 72.230 114.600 72.770 ;
        RECT 115.290 72.550 118.290 72.780 ;
        RECT 114.170 72.170 114.580 72.230 ;
        RECT 117.380 67.040 117.610 68.300 ;
        RECT 118.340 67.050 118.570 68.300 ;
        RECT 119.300 67.080 119.530 68.300 ;
        RECT 117.330 66.510 117.710 67.040 ;
        RECT 118.270 66.520 118.650 67.050 ;
        RECT 117.380 66.300 117.610 66.510 ;
        RECT 118.340 66.300 118.570 66.520 ;
        RECT 119.220 66.460 119.640 67.080 ;
        RECT 119.300 66.300 119.530 66.460 ;
        RECT 116.250 63.250 116.480 63.280 ;
        RECT 117.210 63.250 117.440 63.280 ;
        RECT 116.200 62.620 116.570 63.250 ;
        RECT 117.160 62.620 117.530 63.250 ;
        RECT 118.180 62.750 118.660 63.110 ;
        RECT 116.250 60.280 116.480 62.620 ;
        RECT 117.210 60.280 117.440 62.620 ;
        RECT 121.680 61.650 121.910 61.670 ;
        RECT 121.650 61.340 122.080 61.650 ;
        RECT 121.680 60.670 121.910 61.340 ;
        RECT 119.890 59.970 120.900 59.990 ;
        RECT 119.880 59.650 120.900 59.970 ;
        RECT 119.890 59.610 120.900 59.650 ;
        RECT 114.180 57.300 115.470 58.330 ;
        RECT 105.000 55.640 105.230 55.700 ;
        RECT 104.930 55.360 105.320 55.640 ;
        RECT 105.490 55.370 105.880 55.650 ;
        RECT 105.000 54.700 105.230 55.360 ;
        RECT 95.160 54.120 95.620 54.200 ;
        RECT 95.950 54.120 97.330 54.180 ;
        RECT 95.160 53.720 97.330 54.120 ;
        RECT 95.910 53.710 97.330 53.720 ;
        RECT 95.950 53.700 97.330 53.710 ;
        RECT 26.240 16.160 28.110 16.780 ;
        RECT 15.020 11.690 22.830 12.440 ;
        RECT 3.980 9.100 5.980 11.270 ;
        RECT 20.720 10.920 20.950 11.020 ;
        RECT 20.470 10.010 21.030 10.920 ;
        RECT 23.300 10.840 23.530 11.020 ;
        RECT 23.130 10.170 23.690 10.840 ;
        RECT 25.050 10.780 25.280 14.950 ;
        RECT 23.300 10.020 23.530 10.170 ;
        RECT 24.890 10.030 25.510 10.780 ;
        RECT 27.630 10.730 27.860 14.950 ;
        RECT 25.050 9.950 25.280 10.030 ;
        RECT 27.440 9.980 28.060 10.730 ;
        RECT 30.210 10.710 30.440 14.950 ;
        RECT 32.360 10.960 32.590 19.900 ;
        RECT 27.630 9.950 27.860 9.980 ;
        RECT 30.000 9.960 30.620 10.710 ;
        RECT 32.150 10.190 32.820 10.960 ;
        RECT 34.940 10.950 35.170 19.900 ;
        RECT 30.210 9.950 30.440 9.960 ;
        RECT 32.360 9.900 32.590 10.190 ;
        RECT 34.740 10.180 35.410 10.950 ;
        RECT 37.520 10.850 37.750 19.900 ;
        RECT 34.940 9.900 35.170 10.180 ;
        RECT 37.280 10.080 37.950 10.850 ;
        RECT 99.120 10.090 99.350 16.090 ;
        RECT 102.360 10.090 102.590 16.090 ;
        RECT 104.620 12.230 104.850 16.140 ;
        RECT 106.200 12.230 106.430 16.140 ;
        RECT 107.780 12.230 108.010 16.140 ;
        RECT 109.360 12.230 109.590 16.140 ;
        RECT 37.520 9.900 37.750 10.080 ;
        RECT 21.250 9.180 23.020 9.430 ;
        RECT 26.820 9.180 28.130 9.300 ;
        RECT 21.250 9.130 28.130 9.180 ;
        RECT 34.020 9.130 35.560 9.270 ;
        RECT 39.540 9.130 40.540 9.230 ;
        RECT 20.000 9.100 43.720 9.130 ;
        RECT 3.980 7.160 43.720 9.100 ;
        RECT 98.360 7.270 111.920 8.900 ;
        RECT 3.980 7.130 35.790 7.160 ;
        RECT 3.980 6.700 5.980 7.130 ;
        RECT 3.980 6.600 5.990 6.700 ;
        RECT 99.820 6.600 101.340 7.270 ;
        RECT 3.980 6.090 101.340 6.600 ;
        RECT 4.000 5.080 101.340 6.090 ;
        RECT 4.000 5.040 5.990 5.080 ;
      LAYER met2 ;
        RECT 114.200 72.180 114.550 72.820 ;
        RECT 119.270 67.100 119.590 67.130 ;
        RECT 117.370 66.690 119.590 67.100 ;
        RECT 117.370 66.480 119.630 66.690 ;
        RECT 117.380 66.400 117.680 66.480 ;
        RECT 118.320 66.470 118.600 66.480 ;
        RECT 119.270 66.450 119.620 66.480 ;
        RECT 119.270 66.410 119.590 66.450 ;
        RECT 116.250 63.150 116.520 63.300 ;
        RECT 117.210 63.150 117.480 63.300 ;
        RECT 118.230 63.150 118.610 63.160 ;
        RECT 116.190 62.720 118.660 63.150 ;
        RECT 116.250 62.570 116.520 62.720 ;
        RECT 117.190 62.670 117.490 62.720 ;
        RECT 118.230 62.700 118.610 62.720 ;
        RECT 117.210 62.570 117.480 62.670 ;
        RECT 121.700 61.290 122.030 61.700 ;
        RECT 121.710 61.280 122.000 61.290 ;
        RECT 119.930 59.600 120.820 60.020 ;
        RECT 114.330 57.250 115.420 58.380 ;
        RECT 104.980 55.300 105.300 55.780 ;
        RECT 105.540 55.330 105.890 55.730 ;
        RECT 105.540 55.320 105.830 55.330 ;
        RECT 95.960 53.660 96.330 54.150 ;
        RECT 26.300 16.750 28.050 16.800 ;
        RECT 24.700 16.190 28.050 16.750 ;
        RECT 4.030 6.750 5.930 11.320 ;
        RECT 20.520 10.900 20.980 10.970 ;
        RECT 20.520 10.760 23.690 10.900 ;
        RECT 24.700 10.760 25.490 16.190 ;
        RECT 26.300 16.140 28.050 16.190 ;
        RECT 32.200 10.840 32.770 11.010 ;
        RECT 29.640 10.810 32.980 10.840 ;
        RECT 34.790 10.810 35.360 11.000 ;
        RECT 37.330 10.810 37.900 10.900 ;
        RECT 20.520 10.630 25.490 10.760 ;
        RECT 27.490 10.630 28.010 10.780 ;
        RECT 29.640 10.630 37.900 10.810 ;
        RECT 20.520 10.230 37.900 10.630 ;
        RECT 20.520 10.160 32.980 10.230 ;
        RECT 20.520 10.090 23.690 10.160 ;
        RECT 20.520 9.960 20.980 10.090 ;
        RECT 21.810 9.450 22.370 10.090 ;
        RECT 24.940 10.050 32.980 10.160 ;
        RECT 24.940 10.020 30.570 10.050 ;
        RECT 24.940 9.980 25.460 10.020 ;
        RECT 27.090 9.930 28.010 10.020 ;
        RECT 21.310 8.910 22.960 9.450 ;
        RECT 27.090 9.320 27.930 9.930 ;
        RECT 30.050 9.910 30.570 10.020 ;
        RECT 26.880 8.730 28.070 9.320 ;
        RECT 34.690 9.290 35.430 10.230 ;
        RECT 37.330 10.030 37.900 10.230 ;
        RECT 34.080 8.780 35.500 9.290 ;
        RECT 4.030 6.040 5.940 6.750 ;
        RECT 4.050 4.990 5.940 6.040 ;
      LAYER met3 ;
        RECT 110.060 72.960 112.030 73.520 ;
        RECT 110.060 71.980 114.650 72.960 ;
        RECT 104.930 55.750 105.350 55.755 ;
        RECT 110.060 55.750 112.030 71.980 ;
        RECT 119.280 67.180 119.840 67.370 ;
        RECT 119.230 67.080 119.840 67.180 ;
        RECT 119.220 67.040 119.840 67.080 ;
        RECT 119.220 66.670 119.800 67.040 ;
        RECT 119.220 66.220 119.830 66.670 ;
        RECT 114.280 58.320 115.470 58.355 ;
        RECT 114.080 58.110 115.490 58.320 ;
        RECT 117.130 58.110 117.590 63.270 ;
        RECT 119.220 60.000 119.660 66.220 ;
        RECT 121.690 61.635 122.150 61.650 ;
        RECT 121.660 61.305 122.150 61.635 ;
        RECT 121.690 61.070 122.150 61.305 ;
        RECT 119.220 59.995 120.320 60.000 ;
        RECT 119.220 59.625 120.870 59.995 ;
        RECT 119.220 59.330 120.620 59.625 ;
        RECT 119.220 58.110 119.660 59.330 ;
        RECT 121.810 58.110 122.150 61.070 ;
        RECT 114.080 58.010 120.700 58.110 ;
        RECT 121.510 58.010 122.240 58.110 ;
        RECT 114.080 57.360 122.240 58.010 ;
        RECT 114.080 55.750 115.490 57.360 ;
        RECT 119.220 57.230 119.660 57.360 ;
        RECT 120.320 57.340 121.920 57.360 ;
        RECT 3.970 53.560 5.990 55.590 ;
        RECT 104.930 55.350 115.620 55.750 ;
        RECT 104.930 55.325 105.350 55.350 ;
        RECT 95.800 53.560 96.380 54.170 ;
        RECT 110.060 53.560 112.030 55.350 ;
        RECT 114.080 53.560 115.490 55.350 ;
        RECT 3.970 52.550 115.770 53.560 ;
        RECT 3.970 50.710 5.990 52.550 ;
        RECT 97.760 52.540 99.910 52.550 ;
        RECT 110.060 52.530 112.030 52.550 ;
        RECT 114.080 52.440 115.490 52.550 ;
        RECT 3.980 6.725 5.980 11.295 ;
        RECT 3.980 6.065 5.990 6.725 ;
        RECT 4.000 5.015 5.990 6.065 ;
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 124.640 90.560 138.610 91.990 ;
        RECT 124.640 86.910 126.070 90.560 ;
      LAYER pwell ;
        RECT 126.130 87.020 137.130 90.510 ;
      LAYER nwell ;
        RECT 137.180 86.910 138.610 90.560 ;
        RECT 124.640 85.480 138.610 86.910 ;
        RECT 101.710 74.680 108.670 78.870 ;
        RECT 112.060 73.950 115.650 85.140 ;
      LAYER pwell ;
        RECT 132.085 81.055 135.055 81.485 ;
        RECT 132.085 74.975 132.515 81.055 ;
        RECT 134.625 74.975 135.055 81.055 ;
        RECT 132.085 74.545 135.055 74.975 ;
      LAYER nwell ;
        RECT 101.830 69.120 108.790 73.310 ;
        RECT 102.090 57.660 108.560 67.850 ;
      LAYER pwell ;
        RECT 124.810 64.885 125.740 65.795 ;
        RECT 125.955 64.970 126.385 65.755 ;
        RECT 128.825 65.010 129.255 65.795 ;
        RECT 129.340 64.925 131.250 65.605 ;
        RECT 124.810 64.865 124.915 64.885 ;
        RECT 124.745 64.695 124.915 64.865 ;
        RECT 129.415 64.735 129.585 64.925 ;
        RECT 96.160 54.045 97.090 54.955 ;
        RECT 96.160 54.025 96.265 54.045 ;
        RECT 96.095 53.855 96.265 54.025 ;
      LAYER li1 ;
        RECT 124.925 91.535 138.325 91.705 ;
        RECT 124.925 85.935 125.095 91.535 ;
        RECT 126.260 90.210 137.000 90.380 ;
        RECT 126.260 87.320 126.430 90.210 ;
        RECT 127.110 89.640 136.150 89.810 ;
        RECT 127.110 89.160 136.150 89.330 ;
        RECT 127.110 88.680 136.150 88.850 ;
        RECT 127.110 88.200 136.150 88.370 ;
        RECT 127.110 87.720 136.150 87.890 ;
        RECT 136.830 87.320 137.000 90.210 ;
        RECT 126.260 87.150 137.000 87.320 ;
        RECT 134.010 86.230 135.360 87.150 ;
        RECT 138.155 85.935 138.325 91.535 ;
        RECT 124.925 85.765 138.325 85.935 ;
        RECT 112.240 84.790 115.470 84.960 ;
        RECT 102.590 83.470 107.590 83.640 ;
        RECT 102.360 81.215 102.530 83.255 ;
        RECT 102.590 80.830 107.590 81.000 ;
        RECT 98.900 77.670 100.310 79.830 ;
        RECT 101.890 78.520 108.490 78.690 ;
        RECT 101.890 75.030 102.060 78.520 ;
        RECT 102.690 78.010 107.690 78.180 ;
        RECT 102.460 75.755 102.630 77.795 ;
        RECT 107.750 76.990 107.920 77.795 ;
        RECT 108.320 76.990 108.490 78.520 ;
        RECT 107.750 76.620 108.490 76.990 ;
        RECT 107.750 75.755 107.920 76.620 ;
        RECT 102.690 75.370 107.690 75.540 ;
        RECT 108.320 75.030 108.490 76.620 ;
        RECT 101.890 74.860 108.490 75.030 ;
        RECT 112.240 74.300 112.410 84.790 ;
        RECT 112.810 75.025 112.980 84.065 ;
        RECT 113.290 75.025 113.460 84.065 ;
        RECT 113.770 75.025 113.940 84.065 ;
        RECT 114.250 75.025 114.420 84.065 ;
        RECT 114.730 75.025 114.900 84.065 ;
        RECT 115.300 76.130 115.470 84.790 ;
        RECT 132.215 81.185 134.925 81.355 ;
        RECT 124.260 80.120 124.590 80.290 ;
        RECT 125.220 80.120 125.550 80.290 ;
        RECT 123.780 77.480 124.110 77.650 ;
        RECT 124.740 77.480 125.070 77.650 ;
        RECT 125.700 77.480 126.030 77.650 ;
        RECT 115.300 75.670 115.550 76.130 ;
        RECT 115.300 74.300 115.470 75.670 ;
        RECT 132.215 74.845 132.385 81.185 ;
        RECT 132.865 75.325 134.275 77.485 ;
        RECT 134.755 75.840 134.925 81.185 ;
        RECT 134.720 75.130 148.020 75.840 ;
        RECT 134.755 74.845 134.925 75.130 ;
        RECT 132.215 74.675 134.925 74.845 ;
        RECT 112.240 74.130 115.470 74.300 ;
        RECT 102.010 72.960 108.610 73.130 ;
        RECT 102.010 69.470 102.180 72.960 ;
        RECT 102.810 72.450 107.810 72.620 ;
        RECT 102.580 70.195 102.750 72.235 ;
        RECT 107.870 71.420 108.040 72.235 ;
        RECT 108.440 71.420 108.610 72.960 ;
        RECT 114.930 72.205 115.100 72.535 ;
        RECT 118.480 72.205 118.650 72.535 ;
        RECT 115.270 71.990 118.310 72.160 ;
        RECT 121.230 71.420 146.230 71.590 ;
        RECT 107.870 71.050 108.610 71.420 ;
        RECT 107.870 70.195 108.040 71.050 ;
        RECT 102.810 69.810 107.810 69.980 ;
        RECT 108.440 69.470 108.610 71.050 ;
        RECT 121.230 69.780 146.230 69.950 ;
        RECT 102.010 69.300 108.610 69.470 ;
        RECT 102.270 67.500 108.380 67.670 ;
        RECT 97.900 64.980 99.310 67.140 ;
        RECT 97.900 61.760 99.310 63.920 ;
        RECT 102.270 60.530 102.440 67.500 ;
        RECT 106.380 67.160 106.670 67.200 ;
        RECT 103.480 66.990 103.810 67.160 ;
        RECT 104.440 66.990 104.770 67.160 ;
        RECT 105.400 66.990 105.730 67.160 ;
        RECT 106.360 66.990 106.690 67.160 ;
        RECT 107.320 66.990 107.650 67.160 ;
        RECT 106.380 66.960 106.670 66.990 ;
        RECT 102.020 59.470 102.570 60.530 ;
        RECT 102.270 58.010 102.440 59.470 ;
        RECT 103.320 58.735 103.490 66.775 ;
        RECT 104.280 58.735 104.450 66.775 ;
        RECT 105.240 58.735 105.410 66.775 ;
        RECT 106.200 58.735 106.370 66.775 ;
        RECT 107.160 58.735 107.330 66.775 ;
        RECT 106.860 58.520 107.150 58.560 ;
        RECT 103.000 58.350 103.330 58.520 ;
        RECT 103.960 58.350 104.290 58.520 ;
        RECT 104.920 58.350 105.250 58.520 ;
        RECT 105.880 58.350 106.210 58.520 ;
        RECT 106.840 58.350 107.170 58.520 ;
        RECT 106.860 58.320 107.150 58.350 ;
        RECT 108.210 58.010 108.380 67.500 ;
        RECT 114.700 66.025 114.870 69.065 ;
        RECT 116.930 66.280 117.100 68.320 ;
        RECT 117.890 66.280 118.060 68.320 ;
        RECT 118.850 66.280 119.020 68.320 ;
        RECT 125.320 66.265 125.650 67.245 ;
        RECT 129.870 66.955 130.135 67.285 ;
        RECT 129.400 66.775 129.580 66.780 ;
        RECT 124.920 66.070 125.250 66.095 ;
        RECT 124.860 65.860 125.250 66.070 ;
        RECT 124.920 65.855 125.250 65.860 ;
        RECT 124.920 64.865 125.150 65.685 ;
        RECT 125.420 65.665 125.650 66.265 ;
        RECT 129.355 66.005 129.700 66.775 ;
        RECT 129.870 65.770 130.040 66.955 ;
        RECT 130.230 66.435 130.540 66.460 ;
        RECT 130.210 65.900 130.540 66.435 ;
        RECT 125.320 65.035 125.650 65.665 ;
        RECT 129.455 65.730 130.040 65.770 ;
        RECT 130.720 65.730 131.050 66.255 ;
        RECT 126.025 64.865 126.315 65.590 ;
        RECT 128.895 64.905 129.185 65.630 ;
        RECT 129.455 65.515 131.050 65.730 ;
        RECT 129.455 65.100 129.760 65.515 ;
        RECT 130.220 64.905 130.660 65.345 ;
        RECT 147.510 65.170 147.990 75.130 ;
        RECT 132.340 64.910 148.020 65.170 ;
        RECT 131.530 64.905 148.020 64.910 ;
        RECT 124.600 64.695 126.400 64.865 ;
        RECT 128.810 64.735 148.020 64.905 ;
        RECT 131.530 64.730 148.020 64.735 ;
        RECT 116.440 63.470 116.770 63.640 ;
        RECT 117.400 63.470 117.730 63.640 ;
        RECT 112.730 62.820 113.730 62.990 ;
        RECT 112.500 61.565 112.670 62.605 ;
        RECT 112.730 61.180 113.730 61.350 ;
        RECT 115.800 60.260 115.970 63.300 ;
        RECT 116.760 60.260 116.930 63.300 ;
        RECT 117.720 60.260 117.890 63.300 ;
        RECT 125.550 63.220 126.550 63.390 ;
        RECT 126.840 63.220 127.840 63.390 ;
        RECT 128.130 63.220 129.130 63.390 ;
        RECT 129.420 63.220 130.420 63.390 ;
        RECT 130.710 63.220 131.710 63.390 ;
        RECT 132.000 63.220 133.000 63.390 ;
        RECT 133.290 63.220 134.290 63.390 ;
        RECT 134.580 63.220 135.580 63.390 ;
        RECT 135.870 63.220 136.870 63.390 ;
        RECT 137.160 63.220 138.160 63.390 ;
        RECT 120.650 61.860 121.650 62.030 ;
        RECT 120.420 60.650 120.590 61.690 ;
        RECT 120.650 60.310 121.650 60.480 ;
        RECT 115.960 59.920 116.290 60.090 ;
        RECT 116.920 59.920 117.250 60.090 ;
        RECT 116.940 59.850 117.230 59.920 ;
        RECT 102.270 57.840 108.380 58.010 ;
        RECT 96.670 55.425 97.000 56.405 ;
        RECT 104.730 55.890 105.060 56.060 ;
        RECT 96.270 55.220 96.600 55.255 ;
        RECT 96.250 55.030 96.600 55.220 ;
        RECT 96.270 55.015 96.600 55.030 ;
        RECT 96.770 55.240 97.000 55.425 ;
        RECT 96.770 55.040 97.240 55.240 ;
        RECT 96.770 54.825 97.000 55.040 ;
        RECT 125.320 54.965 125.490 63.005 ;
        RECT 127.900 54.965 128.070 63.005 ;
        RECT 130.480 54.965 130.650 63.005 ;
        RECT 133.060 54.965 133.230 63.005 ;
        RECT 135.640 54.965 135.810 63.005 ;
        RECT 138.220 54.965 138.390 63.005 ;
        RECT 96.670 54.195 97.000 54.825 ;
        RECT 125.550 54.580 126.550 54.750 ;
        RECT 126.840 54.580 127.840 54.750 ;
        RECT 128.130 54.580 129.130 54.750 ;
        RECT 129.420 54.580 130.420 54.750 ;
        RECT 130.710 54.580 131.710 54.750 ;
        RECT 132.000 54.580 133.000 54.750 ;
        RECT 133.290 54.580 134.290 54.750 ;
        RECT 134.580 54.580 135.580 54.750 ;
        RECT 135.870 54.580 136.870 54.750 ;
        RECT 137.160 54.580 138.160 54.750 ;
        RECT 104.730 54.340 105.060 54.510 ;
        RECT 32.775 37.790 33.105 37.960 ;
        RECT 33.365 37.790 33.695 37.960 ;
        RECT 33.955 37.790 34.285 37.960 ;
        RECT 34.545 37.790 34.875 37.960 ;
        RECT 36.805 37.790 37.135 37.960 ;
        RECT 37.395 37.790 37.725 37.960 ;
        RECT 37.985 37.790 38.315 37.960 ;
        RECT 38.575 37.790 38.905 37.960 ;
        RECT 41.275 37.790 41.605 37.960 ;
        RECT 42.255 37.790 42.585 37.960 ;
        RECT 16.890 33.890 17.240 36.050 ;
        RECT 18.900 33.890 19.250 36.050 ;
        RECT 20.900 33.890 21.250 36.050 ;
        RECT 22.910 33.890 23.260 36.050 ;
        RECT 25.220 17.410 25.390 32.450 ;
        RECT 25.810 17.410 25.980 32.450 ;
        RECT 26.400 17.410 26.570 32.450 ;
        RECT 28.070 17.410 28.240 32.450 ;
        RECT 28.660 17.410 28.830 32.450 ;
        RECT 29.250 17.410 29.420 32.450 ;
        RECT 33.150 22.535 33.320 37.575 ;
        RECT 34.330 22.535 34.500 37.575 ;
        RECT 37.180 22.535 37.350 37.575 ;
        RECT 38.360 22.535 38.530 37.575 ;
        RECT 99.365 25.905 99.865 26.075 ;
        RECT 101.780 25.920 102.280 26.090 ;
        RECT 99.925 23.650 100.095 25.690 ;
        RECT 101.550 23.665 101.720 25.705 ;
        RECT 99.365 23.265 99.865 23.435 ;
        RECT 101.780 23.280 102.280 23.450 ;
        RECT 32.775 22.150 33.105 22.320 ;
        RECT 33.365 22.150 33.695 22.320 ;
        RECT 33.955 22.150 34.285 22.320 ;
        RECT 34.545 22.150 34.875 22.320 ;
        RECT 36.805 22.150 37.135 22.320 ;
        RECT 37.395 22.150 37.725 22.320 ;
        RECT 37.985 22.150 38.315 22.320 ;
        RECT 38.575 22.150 38.905 22.320 ;
        RECT 32.620 20.090 33.620 20.260 ;
        RECT 33.910 20.090 34.910 20.260 ;
        RECT 35.200 20.090 36.200 20.260 ;
        RECT 36.490 20.090 37.490 20.260 ;
        RECT 99.105 18.350 99.275 21.390 ;
        RECT 99.895 18.350 100.065 21.390 ;
        RECT 101.560 18.350 101.730 21.390 ;
        RECT 102.350 18.350 102.520 21.390 ;
        RECT 105.840 20.635 106.340 20.805 ;
        RECT 106.630 20.635 107.130 20.805 ;
        RECT 107.420 20.635 107.920 20.805 ;
        RECT 108.210 20.635 108.710 20.805 ;
        RECT 109.000 20.635 109.500 20.805 ;
        RECT 105.310 18.770 105.480 18.850 ;
        RECT 116.280 18.770 116.450 18.850 ;
        RECT 105.310 18.600 107.295 18.770 ;
        RECT 114.465 18.600 116.450 18.770 ;
        RECT 105.310 18.520 105.480 18.600 ;
        RECT 116.280 18.520 116.450 18.600 ;
        RECT 40.785 18.150 41.115 18.320 ;
        RECT 41.765 18.150 42.095 18.320 ;
        RECT 104.880 16.330 105.380 16.500 ;
        RECT 105.670 16.330 106.170 16.500 ;
        RECT 106.460 16.330 106.960 16.500 ;
        RECT 107.250 16.330 107.750 16.500 ;
        RECT 108.040 16.330 108.540 16.500 ;
        RECT 108.830 16.330 109.330 16.500 ;
        RECT 25.310 15.140 26.310 15.310 ;
        RECT 26.600 15.140 27.600 15.310 ;
        RECT 27.890 15.140 28.890 15.310 ;
        RECT 29.180 15.140 30.180 15.310 ;
        RECT 14.890 12.890 15.240 15.050 ;
        RECT 16.890 12.890 17.240 15.050 ;
        RECT 18.900 12.890 19.250 15.050 ;
        RECT 20.900 12.890 21.250 15.050 ;
        RECT 22.910 12.890 23.260 15.050 ;
        RECT 20.980 11.210 21.980 11.380 ;
        RECT 22.270 11.210 23.270 11.380 ;
        RECT 22.040 10.000 22.210 11.040 ;
        RECT 26.370 9.930 26.540 14.970 ;
        RECT 28.950 9.930 29.120 14.970 ;
        RECT 39.850 13.580 40.540 15.740 ;
        RECT 20.980 9.660 21.980 9.830 ;
        RECT 22.270 9.660 23.270 9.830 ;
        RECT 25.310 9.590 26.310 9.760 ;
        RECT 26.600 9.590 27.600 9.760 ;
        RECT 27.890 9.590 28.890 9.760 ;
        RECT 29.180 9.590 30.180 9.760 ;
        RECT 32.620 9.540 33.620 9.710 ;
        RECT 33.910 9.540 34.910 9.710 ;
        RECT 35.200 9.540 36.200 9.710 ;
        RECT 36.490 9.540 37.490 9.710 ;
        RECT 39.660 9.500 40.850 12.130 ;
        RECT 99.940 10.070 100.110 16.110 ;
        RECT 101.600 10.070 101.770 16.110 ;
        RECT 96.120 7.590 96.810 9.750 ;
        RECT 99.380 9.730 99.880 9.900 ;
        RECT 101.830 9.730 102.330 9.900 ;
      LAYER met1 ;
        RECT 128.230 89.840 132.600 89.880 ;
        RECT 127.130 89.610 136.130 89.840 ;
        RECT 133.430 89.360 135.810 89.380 ;
        RECT 127.130 89.130 136.130 89.360 ;
        RECT 133.430 89.110 135.810 89.130 ;
        RECT 128.250 88.880 132.620 88.910 ;
        RECT 127.130 88.650 136.130 88.880 ;
        RECT 133.390 88.400 135.770 88.440 ;
        RECT 127.130 88.170 136.130 88.400 ;
        RECT 127.130 87.690 136.130 87.920 ;
        RECT 128.300 87.650 132.670 87.690 ;
        RECT 119.430 86.630 119.710 86.730 ;
        RECT 133.950 86.630 135.420 87.350 ;
        RECT 119.430 86.200 135.420 86.630 ;
        RECT 119.430 86.020 135.300 86.200 ;
        RECT 102.530 83.750 107.620 83.820 ;
        RECT 102.230 83.380 107.620 83.750 ;
        RECT 102.230 83.230 102.560 83.380 ;
        RECT 102.230 81.240 102.640 83.230 ;
        RECT 112.780 81.460 113.010 84.045 ;
        RECT 102.230 81.090 102.560 81.240 ;
        RECT 102.230 80.650 107.820 81.090 ;
        RECT 112.690 80.680 113.050 81.460 ;
        RECT 98.940 79.750 100.330 79.880 ;
        RECT 98.780 77.810 100.330 79.750 ;
        RECT 104.240 79.800 105.490 80.650 ;
        RECT 108.970 79.800 109.460 79.830 ;
        RECT 104.240 79.300 109.500 79.800 ;
        RECT 102.360 78.300 102.770 78.330 ;
        RECT 102.350 77.920 107.690 78.300 ;
        RECT 98.780 77.700 100.260 77.810 ;
        RECT 96.540 75.160 97.680 75.240 ;
        RECT 98.780 75.160 100.250 77.700 ;
        RECT 102.360 77.560 102.770 77.920 ;
        RECT 102.340 76.350 102.770 77.560 ;
        RECT 107.720 77.240 107.950 77.775 ;
        RECT 108.970 77.240 109.460 79.300 ;
        RECT 102.360 75.620 102.770 76.350 ;
        RECT 107.600 76.330 109.700 77.240 ;
        RECT 107.680 76.320 109.700 76.330 ;
        RECT 107.720 75.775 107.950 76.320 ;
        RECT 108.970 76.300 109.460 76.320 ;
        RECT 104.560 75.620 105.540 75.710 ;
        RECT 102.360 75.300 107.700 75.620 ;
        RECT 102.360 75.170 102.770 75.300 ;
        RECT 96.540 74.100 100.250 75.160 ;
        RECT 104.560 74.990 105.540 75.300 ;
        RECT 112.780 75.045 113.010 80.680 ;
        RECT 113.260 76.290 113.490 84.045 ;
        RECT 113.740 81.450 113.970 84.045 ;
        RECT 113.700 80.670 114.060 81.450 ;
        RECT 113.190 75.510 113.550 76.290 ;
        RECT 113.260 75.045 113.490 75.510 ;
        RECT 113.740 75.045 113.970 80.670 ;
        RECT 114.220 76.260 114.450 84.045 ;
        RECT 114.700 81.480 114.930 84.045 ;
        RECT 114.640 80.700 115.000 81.480 ;
        RECT 114.180 75.480 114.540 76.260 ;
        RECT 114.220 75.045 114.450 75.480 ;
        RECT 114.700 75.045 114.930 80.700 ;
        RECT 115.270 76.170 115.580 76.190 ;
        RECT 115.250 75.700 115.630 76.170 ;
        RECT 115.270 75.610 115.580 75.700 ;
        RECT 104.580 74.360 105.530 74.990 ;
        RECT 109.120 74.360 109.670 74.370 ;
        RECT 96.540 69.970 97.680 74.100 ;
        RECT 98.780 74.090 100.250 74.100 ;
        RECT 104.540 73.930 109.670 74.360 ;
        RECT 105.120 73.920 109.670 73.930 ;
        RECT 102.520 72.710 102.840 72.720 ;
        RECT 102.520 72.370 107.810 72.710 ;
        RECT 102.520 72.210 102.840 72.370 ;
        RECT 102.450 70.220 102.860 72.210 ;
        RECT 107.750 71.840 108.300 72.230 ;
        RECT 107.750 71.600 108.280 71.840 ;
        RECT 109.120 71.600 109.670 73.920 ;
        RECT 114.780 72.780 115.090 73.030 ;
        RECT 114.780 72.390 115.150 72.780 ;
        RECT 118.450 72.390 118.700 72.820 ;
        RECT 114.780 72.380 118.820 72.390 ;
        RECT 119.430 72.380 119.710 86.020 ;
        RECT 121.570 83.870 122.500 83.890 ;
        RECT 120.970 82.790 123.000 83.870 ;
        RECT 121.570 80.410 122.500 82.790 ;
        RECT 121.570 80.400 124.130 80.410 ;
        RECT 121.570 80.040 126.230 80.400 ;
        RECT 121.570 80.030 124.130 80.040 ;
        RECT 121.570 77.720 122.500 80.030 ;
        RECT 121.570 77.710 124.740 77.720 ;
        RECT 121.570 77.350 126.190 77.710 ;
        RECT 132.915 77.430 134.225 77.460 ;
        RECT 121.570 77.290 124.740 77.350 ;
        RECT 122.260 77.270 124.740 77.290 ;
        RECT 132.790 75.400 134.300 77.430 ;
        RECT 132.915 75.355 134.225 75.400 ;
        RECT 114.790 72.150 119.920 72.380 ;
        RECT 114.790 72.140 118.820 72.150 ;
        RECT 114.850 72.110 118.820 72.140 ;
        RECT 119.430 72.130 119.710 72.150 ;
        RECT 115.290 71.960 118.290 72.110 ;
        RECT 107.750 70.950 109.670 71.600 ;
        RECT 121.250 71.390 146.210 71.620 ;
        RECT 107.750 70.840 108.280 70.950 ;
        RECT 107.730 70.250 108.260 70.840 ;
        RECT 102.520 70.020 102.840 70.220 ;
        RECT 107.840 70.215 108.070 70.250 ;
        RECT 100.610 70.010 103.080 70.020 ;
        RECT 100.610 69.980 107.790 70.010 ;
        RECT 96.540 68.980 99.310 69.970 ;
        RECT 96.580 68.970 99.310 68.980 ;
        RECT 97.990 67.130 99.310 68.970 ;
        RECT 100.580 69.780 107.790 69.980 ;
        RECT 121.250 69.960 146.210 69.980 ;
        RECT 100.580 69.730 107.770 69.780 ;
        RECT 120.990 69.750 146.210 69.960 ;
        RECT 100.580 69.650 103.080 69.730 ;
        RECT 97.890 64.960 99.370 67.130 ;
        RECT 97.990 64.950 99.310 64.960 ;
        RECT 97.950 63.780 99.260 63.895 ;
        RECT 95.200 63.350 97.530 63.360 ;
        RECT 97.890 63.350 99.370 63.780 ;
        RECT 92.680 63.330 94.050 63.340 ;
        RECT 95.200 63.330 99.430 63.350 ;
        RECT 92.680 61.920 99.430 63.330 ;
        RECT 92.680 61.890 95.360 61.920 ;
        RECT 97.100 61.890 99.430 61.920 ;
        RECT 92.680 55.280 94.050 61.890 ;
        RECT 97.890 61.610 99.370 61.890 ;
        RECT 100.580 60.550 101.480 69.650 ;
        RECT 114.670 68.530 114.900 69.045 ;
        RECT 114.390 67.740 114.960 68.530 ;
        RECT 116.900 68.230 117.130 68.300 ;
        RECT 107.310 67.310 109.650 67.480 ;
        RECT 103.470 66.900 109.650 67.310 ;
        RECT 103.290 61.170 103.520 66.755 ;
        RECT 104.250 61.220 104.480 66.755 ;
        RECT 100.610 60.510 101.620 60.550 ;
        RECT 101.990 60.510 102.600 60.590 ;
        RECT 103.200 60.510 103.590 61.170 ;
        RECT 100.610 59.590 102.600 60.510 ;
        RECT 103.290 59.590 103.520 60.510 ;
        RECT 100.610 59.570 101.620 59.590 ;
        RECT 101.990 59.410 102.600 59.590 ;
        RECT 103.200 58.890 103.590 59.590 ;
        RECT 104.170 58.940 104.560 61.220 ;
        RECT 105.210 61.210 105.440 66.755 ;
        RECT 103.290 58.755 103.520 58.890 ;
        RECT 104.250 58.755 104.480 58.940 ;
        RECT 105.130 58.930 105.520 61.210 ;
        RECT 106.170 61.140 106.400 66.755 ;
        RECT 107.130 61.140 107.360 66.755 ;
        RECT 105.210 58.755 105.440 58.930 ;
        RECT 106.090 58.860 106.480 61.140 ;
        RECT 107.050 58.860 107.440 61.140 ;
        RECT 106.170 58.755 106.400 58.860 ;
        RECT 107.130 58.755 107.360 58.860 ;
        RECT 109.240 58.610 109.650 66.900 ;
        RECT 114.670 66.045 114.900 67.740 ;
        RECT 116.800 67.700 117.180 68.230 ;
        RECT 117.860 68.220 118.090 68.300 ;
        RECT 116.900 66.300 117.130 67.700 ;
        RECT 117.760 67.690 118.140 68.220 ;
        RECT 118.820 68.210 119.050 68.300 ;
        RECT 117.860 66.300 118.090 67.690 ;
        RECT 118.770 67.680 119.150 68.210 ;
        RECT 120.990 68.070 122.450 69.750 ;
        RECT 118.820 66.300 119.050 67.680 ;
        RECT 120.980 67.340 122.450 68.070 ;
        RECT 120.990 67.290 122.450 67.340 ;
        RECT 121.010 67.240 121.990 67.290 ;
        RECT 121.030 66.230 121.990 67.240 ;
        RECT 129.370 66.830 129.610 66.840 ;
        RECT 129.310 66.490 129.710 66.830 ;
        RECT 125.420 66.430 126.560 66.450 ;
        RECT 125.360 66.320 126.560 66.430 ;
        RECT 130.170 66.320 130.600 66.490 ;
        RECT 125.360 66.260 130.600 66.320 ;
        RECT 121.030 66.130 122.280 66.230 ;
        RECT 125.360 66.200 125.950 66.260 ;
        RECT 126.290 66.190 130.600 66.260 ;
        RECT 126.290 66.180 130.560 66.190 ;
        RECT 121.030 66.090 124.290 66.130 ;
        RECT 121.030 65.900 125.200 66.090 ;
        RECT 120.890 65.820 125.200 65.900 ;
        RECT 120.890 65.550 124.290 65.820 ;
        RECT 114.610 64.910 115.430 65.300 ;
        RECT 120.890 65.080 122.420 65.550 ;
        RECT 129.090 65.200 129.840 65.290 ;
        RECT 119.870 64.650 122.570 65.080 ;
        RECT 119.860 64.240 122.570 64.650 ;
        RECT 124.500 65.020 125.160 65.140 ;
        RECT 128.930 65.060 129.840 65.200 ;
        RECT 124.500 64.640 126.400 65.020 ;
        RECT 124.570 64.540 126.400 64.640 ;
        RECT 128.810 64.580 131.570 65.060 ;
        RECT 111.530 63.850 117.980 63.860 ;
        RECT 119.860 63.850 120.270 64.240 ;
        RECT 121.950 64.170 122.310 64.240 ;
        RECT 111.530 63.440 120.270 63.850 ;
        RECT 126.980 63.510 137.600 63.560 ;
        RECT 111.530 63.430 119.980 63.440 ;
        RECT 111.530 63.420 117.980 63.430 ;
        RECT 122.980 63.420 137.600 63.510 ;
        RECT 111.540 63.090 112.080 63.420 ;
        RECT 111.540 62.850 113.720 63.090 ;
        RECT 111.550 62.760 113.720 62.850 ;
        RECT 111.550 61.470 112.070 62.760 ;
        RECT 112.470 62.050 112.700 62.585 ;
        RECT 115.770 62.050 116.000 63.280 ;
        RECT 112.320 61.630 112.750 62.050 ;
        RECT 115.650 61.630 116.080 62.050 ;
        RECT 116.730 62.040 116.960 63.280 ;
        RECT 117.690 62.050 117.920 63.280 ;
        RECT 122.980 63.190 138.140 63.420 ;
        RECT 122.980 63.150 137.600 63.190 ;
        RECT 122.980 63.130 123.380 63.150 ;
        RECT 122.740 63.000 123.380 63.130 ;
        RECT 122.740 62.220 123.300 63.000 ;
        RECT 122.710 62.210 123.450 62.220 ;
        RECT 119.600 62.190 123.450 62.210 ;
        RECT 112.470 61.585 112.700 61.630 ;
        RECT 111.550 61.350 112.100 61.470 ;
        RECT 112.750 61.350 113.710 61.380 ;
        RECT 111.550 61.070 113.800 61.350 ;
        RECT 111.560 61.060 113.800 61.070 ;
        RECT 111.560 60.130 112.100 61.060 ;
        RECT 115.770 60.280 116.000 61.630 ;
        RECT 116.640 61.620 117.070 62.040 ;
        RECT 117.620 62.030 118.050 62.050 ;
        RECT 119.550 62.030 123.450 62.190 ;
        RECT 117.620 61.830 123.450 62.030 ;
        RECT 125.290 61.970 125.520 62.985 ;
        RECT 127.870 62.040 128.100 62.985 ;
        RECT 117.620 61.810 121.880 61.830 ;
        RECT 117.620 61.630 120.020 61.810 ;
        RECT 116.730 60.280 116.960 61.620 ;
        RECT 117.690 61.570 120.020 61.630 ;
        RECT 117.690 60.280 117.920 61.570 ;
        RECT 119.550 61.480 120.010 61.570 ;
        RECT 119.610 60.530 119.930 61.480 ;
        RECT 120.390 61.000 120.620 61.670 ;
        RECT 122.710 61.140 123.450 61.830 ;
        RECT 120.330 60.680 120.690 61.000 ;
        RECT 122.720 60.800 123.450 61.140 ;
        RECT 120.390 60.670 120.620 60.680 ;
        RECT 119.530 60.130 121.810 60.530 ;
        RECT 111.560 59.660 118.500 60.130 ;
        RECT 111.560 59.610 112.100 59.660 ;
        RECT 102.940 58.580 106.190 58.610 ;
        RECT 106.600 58.580 109.650 58.610 ;
        RECT 102.940 58.240 109.650 58.580 ;
        RECT 106.080 57.300 106.490 58.240 ;
        RECT 106.640 58.190 109.650 58.240 ;
        RECT 97.800 56.780 106.500 57.300 ;
        RECT 97.800 55.290 98.200 56.780 ;
        RECT 106.080 56.180 106.490 56.780 ;
        RECT 104.630 55.920 106.490 56.180 ;
        RECT 104.630 55.840 106.590 55.920 ;
        RECT 92.640 54.900 96.580 55.280 ;
        RECT 96.960 55.270 98.210 55.290 ;
        RECT 96.900 55.210 98.210 55.270 ;
        RECT 96.900 55.010 98.220 55.210 ;
        RECT 96.980 54.990 98.220 55.010 ;
        RECT 106.180 54.550 106.590 55.840 ;
        RECT 122.710 54.840 123.450 60.800 ;
        RECT 125.120 60.750 125.670 61.970 ;
        RECT 127.730 60.780 128.250 62.040 ;
        RECT 130.450 61.960 130.680 62.985 ;
        RECT 125.290 54.985 125.520 60.750 ;
        RECT 127.870 54.985 128.100 60.780 ;
        RECT 130.310 60.700 130.830 61.960 ;
        RECT 133.030 61.920 133.260 62.985 ;
        RECT 135.610 61.920 135.840 62.985 ;
        RECT 138.190 61.990 138.420 62.985 ;
        RECT 130.450 54.985 130.680 60.700 ;
        RECT 132.900 60.660 133.420 61.920 ;
        RECT 135.460 60.660 135.980 61.920 ;
        RECT 138.020 60.730 138.540 61.990 ;
        RECT 133.030 54.985 133.260 60.660 ;
        RECT 135.610 54.985 135.840 60.660 ;
        RECT 138.190 54.985 138.420 60.730 ;
        RECT 104.530 54.140 106.590 54.550 ;
        RECT 122.530 54.780 137.660 54.840 ;
        RECT 122.530 54.550 138.140 54.780 ;
        RECT 122.530 54.420 137.660 54.550 ;
        RECT 32.850 37.990 39.160 38.080 ;
        RECT 32.795 37.760 39.160 37.990 ;
        RECT 32.850 37.740 39.160 37.760 ;
        RECT 39.700 37.990 40.100 38.050 ;
        RECT 39.700 37.750 42.570 37.990 ;
        RECT 33.020 36.840 33.530 37.740 ;
        RECT 34.290 36.870 34.660 37.740 ;
        RECT 16.940 35.330 17.190 36.020 ;
        RECT 18.950 35.330 19.200 36.020 ;
        RECT 16.940 34.650 19.200 35.330 ;
        RECT 16.940 33.915 17.190 34.650 ;
        RECT 18.950 33.915 19.200 34.650 ;
        RECT 20.950 35.320 21.200 36.020 ;
        RECT 22.960 35.320 23.210 36.020 ;
        RECT 20.950 34.780 23.210 35.320 ;
        RECT 20.950 33.915 21.200 34.780 ;
        RECT 22.960 33.915 23.210 34.780 ;
        RECT 25.190 18.750 25.420 32.430 ;
        RECT 25.780 31.050 26.010 32.430 ;
        RECT 25.690 29.580 26.210 31.050 ;
        RECT 25.040 17.890 25.580 18.750 ;
        RECT 25.190 17.430 25.420 17.890 ;
        RECT 25.780 17.430 26.010 29.580 ;
        RECT 26.370 18.710 26.600 32.430 ;
        RECT 28.040 18.730 28.270 32.430 ;
        RECT 28.630 24.440 28.860 32.430 ;
        RECT 28.500 23.240 29.000 24.440 ;
        RECT 26.210 17.850 26.750 18.710 ;
        RECT 27.910 17.900 28.370 18.730 ;
        RECT 26.370 17.430 26.600 17.850 ;
        RECT 28.040 17.430 28.270 17.900 ;
        RECT 28.630 17.430 28.860 23.240 ;
        RECT 29.220 18.720 29.450 32.430 ;
        RECT 33.120 31.040 33.350 36.840 ;
        RECT 34.300 31.040 34.530 36.870 ;
        RECT 33.040 29.570 33.560 31.040 ;
        RECT 34.210 29.570 34.730 31.040 ;
        RECT 33.120 23.040 33.350 29.570 ;
        RECT 34.300 23.120 34.530 29.570 ;
        RECT 33.090 22.360 33.460 23.040 ;
        RECT 34.260 22.360 34.630 23.120 ;
        RECT 35.590 22.360 36.080 37.740 ;
        RECT 37.150 24.450 37.380 37.555 ;
        RECT 37.020 23.250 37.520 24.450 ;
        RECT 38.330 24.420 38.560 37.555 ;
        RECT 39.700 24.440 40.100 37.750 ;
        RECT 99.385 26.090 99.845 26.105 ;
        RECT 101.800 26.090 102.260 26.120 ;
        RECT 99.350 25.890 102.300 26.090 ;
        RECT 99.385 25.875 100.140 25.890 ;
        RECT 99.900 25.670 100.140 25.875 ;
        RECT 99.895 25.490 100.140 25.670 ;
        RECT 37.150 22.555 37.380 23.250 ;
        RECT 38.190 23.220 38.690 24.420 ;
        RECT 39.640 23.250 40.140 24.440 ;
        RECT 99.895 24.020 100.125 25.490 ;
        RECT 101.520 24.020 101.750 25.685 ;
        RECT 99.895 23.840 100.670 24.020 ;
        RECT 99.895 23.670 100.125 23.840 ;
        RECT 38.330 22.555 38.560 23.220 ;
        RECT 32.740 22.060 39.100 22.360 ;
        RECT 31.140 20.400 31.640 20.480 ;
        RECT 31.140 20.070 37.600 20.400 ;
        RECT 29.120 17.890 29.580 18.720 ;
        RECT 29.220 17.430 29.450 17.890 ;
        RECT 24.100 15.350 24.360 15.450 ;
        RECT 31.140 15.390 31.640 20.070 ;
        RECT 32.640 20.060 33.600 20.070 ;
        RECT 33.930 20.060 34.890 20.070 ;
        RECT 35.220 20.060 36.180 20.070 ;
        RECT 36.510 20.060 37.470 20.070 ;
        RECT 39.700 18.340 40.100 23.250 ;
        RECT 99.385 23.235 99.845 23.465 ;
        RECT 99.075 18.670 99.305 21.370 ;
        RECT 98.480 18.430 99.305 18.670 ;
        RECT 40.805 18.340 41.095 18.350 ;
        RECT 41.785 18.340 42.075 18.350 ;
        RECT 39.640 18.100 42.350 18.340 ;
        RECT 39.700 18.080 40.740 18.100 ;
        RECT 30.130 15.350 31.640 15.390 ;
        RECT 24.100 15.110 31.640 15.350 ;
        RECT 24.100 15.100 30.240 15.110 ;
        RECT 14.940 14.050 15.190 15.025 ;
        RECT 16.940 14.050 17.190 15.025 ;
        RECT 14.940 13.370 17.190 14.050 ;
        RECT 14.940 12.920 15.190 13.370 ;
        RECT 16.940 12.920 17.190 13.370 ;
        RECT 18.950 14.020 19.200 15.025 ;
        RECT 20.950 14.020 21.200 15.025 ;
        RECT 18.950 13.340 21.200 14.020 ;
        RECT 18.950 12.920 19.200 13.340 ;
        RECT 20.950 12.920 21.200 13.340 ;
        RECT 22.960 14.190 23.210 15.025 ;
        RECT 24.100 14.190 24.360 15.100 ;
        RECT 26.340 14.710 26.570 14.950 ;
        RECT 28.920 14.710 29.150 14.950 ;
        RECT 22.960 13.540 24.360 14.190 ;
        RECT 26.140 13.960 26.760 14.710 ;
        RECT 28.730 13.960 29.350 14.710 ;
        RECT 22.960 12.920 23.210 13.540 ;
        RECT 24.100 11.530 24.360 13.540 ;
        RECT 24.100 11.520 24.370 11.530 ;
        RECT 20.980 11.400 21.970 11.520 ;
        RECT 22.290 11.400 24.370 11.520 ;
        RECT 20.980 11.240 24.370 11.400 ;
        RECT 20.980 11.230 23.250 11.240 ;
        RECT 21.000 11.180 23.250 11.230 ;
        RECT 21.920 10.750 22.370 11.180 ;
        RECT 22.010 10.020 22.240 10.750 ;
        RECT 24.100 9.870 24.370 11.240 ;
        RECT 26.340 9.950 26.570 13.960 ;
        RECT 28.920 9.950 29.150 13.960 ;
        RECT 20.980 9.780 24.370 9.870 ;
        RECT 25.330 9.780 26.290 9.790 ;
        RECT 26.620 9.780 27.580 9.790 ;
        RECT 27.910 9.780 28.870 9.790 ;
        RECT 29.200 9.780 30.160 9.790 ;
        RECT 20.980 9.770 30.230 9.780 ;
        RECT 31.140 9.770 31.640 15.110 ;
        RECT 39.730 14.260 40.740 18.080 ;
        RECT 98.480 17.670 98.720 18.430 ;
        RECT 99.075 18.370 99.305 18.430 ;
        RECT 99.865 21.320 100.095 21.370 ;
        RECT 100.460 21.320 100.670 23.840 ;
        RECT 99.865 21.140 100.670 21.320 ;
        RECT 100.980 23.840 101.750 24.020 ;
        RECT 100.980 22.590 101.190 23.840 ;
        RECT 101.520 23.685 101.750 23.840 ;
        RECT 101.800 23.250 102.260 23.480 ;
        RECT 100.980 22.420 104.160 22.590 ;
        RECT 100.980 21.330 101.190 22.420 ;
        RECT 101.530 21.330 101.760 21.370 ;
        RECT 100.980 21.150 101.760 21.330 ;
        RECT 99.865 18.370 100.095 21.140 ;
        RECT 101.530 18.370 101.760 21.150 ;
        RECT 102.320 18.780 102.550 21.370 ;
        RECT 104.000 20.830 104.160 22.420 ;
        RECT 105.860 20.830 106.320 20.835 ;
        RECT 106.650 20.830 107.110 20.835 ;
        RECT 107.440 20.830 107.900 20.835 ;
        RECT 108.230 20.830 108.690 20.835 ;
        RECT 109.020 20.830 109.480 20.835 ;
        RECT 104.000 20.630 109.480 20.830 ;
        RECT 104.000 18.840 104.150 20.630 ;
        RECT 105.860 20.605 106.320 20.630 ;
        RECT 106.650 20.605 107.110 20.630 ;
        RECT 107.440 20.605 107.900 20.630 ;
        RECT 108.230 20.605 108.690 20.630 ;
        RECT 109.020 20.605 109.480 20.630 ;
        RECT 104.000 18.800 105.500 18.840 ;
        RECT 116.200 18.800 116.600 18.890 ;
        RECT 102.320 18.540 103.100 18.780 ;
        RECT 102.320 18.370 102.550 18.540 ;
        RECT 102.910 17.670 103.100 18.540 ;
        RECT 104.000 18.570 107.355 18.800 ;
        RECT 114.405 18.570 116.600 18.800 ;
        RECT 104.000 18.490 105.500 18.570 ;
        RECT 98.480 17.660 103.100 17.670 ;
        RECT 98.480 17.490 103.090 17.660 ;
        RECT 39.900 13.605 40.490 14.260 ;
        RECT 39.630 12.130 40.880 12.190 ;
        RECT 20.980 9.760 31.640 9.770 ;
        RECT 20.980 9.590 37.500 9.760 ;
        RECT 20.980 9.580 23.200 9.590 ;
        RECT 24.100 9.470 37.500 9.590 ;
        RECT 39.610 9.500 40.900 12.130 ;
        RECT 99.910 10.290 100.140 16.090 ;
        RECT 101.550 15.840 101.850 17.490 ;
        RECT 103.400 16.530 103.900 16.540 ;
        RECT 103.400 16.300 109.310 16.530 ;
        RECT 103.400 16.290 103.900 16.300 ;
        RECT 99.900 10.090 100.140 10.290 ;
        RECT 101.570 10.090 101.800 15.840 ;
        RECT 99.900 9.940 100.100 10.090 ;
        RECT 99.400 9.890 102.350 9.940 ;
        RECT 103.400 9.890 103.600 16.290 ;
        RECT 116.200 13.440 116.600 18.570 ;
        RECT 116.200 12.640 149.650 13.440 ;
        RECT 96.170 9.710 96.760 9.725 ;
        RECT 99.400 9.710 103.600 9.890 ;
        RECT 96.110 9.690 103.600 9.710 ;
        RECT 24.100 9.430 24.360 9.470 ;
        RECT 31.140 9.380 31.640 9.470 ;
        RECT 39.630 9.440 40.880 9.500 ;
        RECT 96.110 9.400 99.910 9.690 ;
        RECT 96.110 9.390 98.180 9.400 ;
        RECT 99.400 9.390 99.860 9.400 ;
        RECT 96.170 7.620 96.760 9.390 ;
      LAYER met2 ;
        RECT 128.280 89.570 132.550 89.930 ;
        RECT 129.450 88.960 131.100 89.570 ;
        RECT 133.480 89.060 135.760 89.430 ;
        RECT 128.300 88.600 132.570 88.960 ;
        RECT 129.450 87.960 131.100 88.600 ;
        RECT 134.040 88.490 135.330 89.060 ;
        RECT 133.440 88.120 135.720 88.490 ;
        RECT 128.350 87.600 132.620 87.960 ;
        RECT 129.450 86.930 131.100 87.600 ;
        RECT 134.040 87.370 135.330 88.120 ;
        RECT 129.605 84.030 130.795 86.930 ;
        RECT 134.010 86.180 135.360 87.370 ;
        RECT 134.040 86.130 135.330 86.180 ;
        RECT 121.020 83.900 122.950 83.920 ;
        RECT 129.450 83.900 131.100 84.030 ;
        RECT 102.280 81.190 102.590 83.280 ;
        RECT 116.980 82.840 131.130 83.900 ;
        RECT 116.980 81.760 118.040 82.840 ;
        RECT 121.020 82.740 122.950 82.840 ;
        RECT 112.790 81.510 118.040 81.760 ;
        RECT 112.740 80.700 118.040 81.510 ;
        RECT 112.740 80.630 113.000 80.700 ;
        RECT 113.750 80.620 114.010 80.700 ;
        RECT 114.690 80.650 114.950 80.700 ;
        RECT 98.990 77.760 100.280 79.930 ;
        RECT 102.390 76.300 102.660 77.610 ;
        RECT 107.650 76.280 108.040 77.290 ;
        RECT 108.310 76.410 108.600 77.250 ;
        RECT 113.240 76.280 113.500 76.340 ;
        RECT 114.230 76.280 114.490 76.310 ;
        RECT 113.240 76.270 114.510 76.280 ;
        RECT 115.290 76.270 115.670 76.400 ;
        RECT 113.240 75.520 115.680 76.270 ;
        RECT 113.240 75.460 113.500 75.520 ;
        RECT 114.180 75.510 115.680 75.520 ;
        RECT 114.230 75.430 114.490 75.510 ;
        RECT 132.840 75.350 134.250 77.480 ;
        RECT 102.500 70.170 102.810 72.260 ;
        RECT 116.550 72.020 117.230 72.390 ;
        RECT 107.810 70.790 108.130 71.980 ;
        RECT 108.440 70.910 108.740 71.650 ;
        RECT 107.820 70.740 108.090 70.790 ;
        RECT 96.630 68.920 97.600 70.050 ;
        RECT 114.440 68.300 114.910 68.580 ;
        RECT 114.350 68.260 119.170 68.300 ;
        RECT 114.350 68.040 122.020 68.260 ;
        RECT 114.350 67.770 122.010 68.040 ;
        RECT 114.440 67.690 114.910 67.770 ;
        RECT 116.850 67.650 117.130 67.770 ;
        RECT 117.810 67.640 118.090 67.770 ;
        RECT 118.820 67.660 122.010 67.770 ;
        RECT 118.820 67.630 119.100 67.660 ;
        RECT 121.030 67.380 122.010 67.660 ;
        RECT 121.030 67.240 122.020 67.380 ;
        RECT 97.940 64.910 99.320 67.180 ;
        RECT 129.360 66.840 129.660 66.880 ;
        RECT 127.770 66.480 129.670 66.840 ;
        RECT 127.780 66.330 128.190 66.480 ;
        RECT 129.360 66.440 129.660 66.480 ;
        RECT 114.660 64.860 115.380 65.350 ;
        RECT 124.570 64.590 125.030 65.010 ;
        RECT 97.940 61.560 99.320 63.830 ;
        RECT 127.780 62.090 128.020 66.330 ;
        RECT 129.140 65.280 129.790 65.340 ;
        RECT 129.130 64.720 129.790 65.280 ;
        RECT 129.130 64.690 129.750 64.720 ;
        RECT 112.370 61.940 112.700 62.060 ;
        RECT 115.700 62.050 116.030 62.060 ;
        RECT 117.670 62.050 118.000 62.060 ;
        RECT 127.780 62.050 128.200 62.090 ;
        RECT 115.700 61.940 118.080 62.050 ;
        RECT 125.310 62.020 138.550 62.050 ;
        RECT 125.170 61.950 138.550 62.020 ;
        RECT 124.230 61.940 138.550 61.950 ;
        RECT 112.370 61.550 118.080 61.940 ;
        RECT 124.180 61.930 138.550 61.940 ;
        RECT 112.370 61.540 116.030 61.550 ;
        RECT 112.700 61.440 115.700 61.540 ;
        RECT 116.690 61.530 117.020 61.550 ;
        RECT 117.670 61.540 118.000 61.550 ;
        RECT 103.250 61.080 103.540 61.220 ;
        RECT 104.220 61.080 104.510 61.270 ;
        RECT 105.180 61.080 105.470 61.260 ;
        RECT 106.140 61.080 106.430 61.190 ;
        RECT 107.100 61.080 107.390 61.190 ;
        RECT 103.080 61.010 107.510 61.080 ;
        RECT 101.470 59.500 107.510 61.010 ;
        RECT 120.380 60.990 120.640 61.050 ;
        RECT 124.150 60.990 138.550 61.930 ;
        RECT 120.380 60.740 138.550 60.990 ;
        RECT 120.380 60.630 120.640 60.740 ;
        RECT 124.150 60.730 138.550 60.740 ;
        RECT 124.150 60.720 125.940 60.730 ;
        RECT 124.230 60.710 125.940 60.720 ;
        RECT 125.170 60.700 125.620 60.710 ;
        RECT 130.360 60.650 130.780 60.730 ;
        RECT 132.950 60.610 133.370 60.730 ;
        RECT 135.510 60.610 135.930 60.730 ;
        RECT 138.070 60.680 138.490 60.730 ;
        RECT 103.080 58.910 107.510 59.500 ;
        RECT 103.250 58.840 103.540 58.910 ;
        RECT 104.220 58.890 104.510 58.910 ;
        RECT 105.180 58.880 105.470 58.910 ;
        RECT 106.140 58.810 106.430 58.910 ;
        RECT 107.100 58.810 107.390 58.910 ;
        RECT 25.740 30.680 26.160 31.100 ;
        RECT 33.090 30.680 33.510 31.090 ;
        RECT 34.260 30.680 34.680 31.090 ;
        RECT 25.740 29.910 34.680 30.680 ;
        RECT 25.740 29.530 26.160 29.910 ;
        RECT 33.090 29.520 33.510 29.910 ;
        RECT 34.260 29.520 34.680 29.910 ;
        RECT 28.550 24.110 28.950 24.490 ;
        RECT 37.070 24.110 37.470 24.500 ;
        RECT 38.240 24.110 38.640 24.470 ;
        RECT 39.690 24.110 40.090 24.490 ;
        RECT 28.550 23.480 40.090 24.110 ;
        RECT 28.550 23.190 28.950 23.480 ;
        RECT 37.070 23.200 37.470 23.480 ;
        RECT 38.240 23.170 38.640 23.480 ;
        RECT 39.690 23.200 40.090 23.480 ;
        RECT 25.090 18.510 25.530 18.800 ;
        RECT 26.260 18.510 26.700 18.760 ;
        RECT 27.960 18.510 28.320 18.780 ;
        RECT 29.170 18.510 29.530 18.770 ;
        RECT 25.090 17.980 29.530 18.510 ;
        RECT 25.090 17.840 25.530 17.980 ;
        RECT 26.260 17.800 26.700 17.980 ;
        RECT 27.960 17.850 28.320 17.980 ;
        RECT 28.570 17.840 29.530 17.980 ;
        RECT 26.190 14.610 26.710 14.760 ;
        RECT 28.570 14.610 29.390 17.840 ;
        RECT 26.190 14.560 29.390 14.610 ;
        RECT 26.190 14.040 29.300 14.560 ;
        RECT 26.190 13.910 26.710 14.040 ;
        RECT 28.780 13.910 29.300 14.040 ;
        RECT 149.250 12.640 149.650 13.440 ;
        RECT 39.660 9.450 40.850 12.180 ;
      LAYER met3 ;
        RECT 132.840 77.455 134.360 77.480 ;
        RECT 115.260 76.375 115.730 76.440 ;
        RECT 115.240 75.615 115.730 76.375 ;
        RECT 115.260 74.720 115.730 75.615 ;
        RECT 132.790 75.375 134.360 77.455 ;
        RECT 132.840 74.720 134.360 75.375 ;
        RECT 115.250 73.720 134.550 74.720 ;
        RECT 129.090 65.260 129.750 65.330 ;
        RECT 129.090 65.255 129.850 65.260 ;
        RECT 124.500 65.020 125.160 65.140 ;
        RECT 129.080 65.020 129.850 65.255 ;
        RECT 124.500 64.720 129.850 65.020 ;
        RECT 124.500 64.700 129.830 64.720 ;
        RECT 124.500 64.640 129.750 64.700 ;
        RECT 124.520 64.615 129.750 64.640 ;
        RECT 124.530 64.610 129.750 64.615 ;
        RECT 124.600 64.550 129.730 64.610 ;
        RECT 117.850 13.890 149.710 44.290 ;
        RECT 149.250 12.640 149.650 13.890 ;
        RECT 39.610 9.475 40.900 12.155 ;
      LAYER met4 ;
        RECT 149.210 13.950 149.690 44.230 ;
        RECT 38.770 9.470 41.590 12.450 ;
      LAYER met5 ;
        RECT 38.650 11.660 41.710 12.570 ;
        RECT 44.970 11.660 74.810 39.005 ;
        RECT 38.650 9.790 74.810 11.660 ;
        RECT 38.650 9.350 41.710 9.790 ;
        RECT 44.970 9.165 74.810 9.790 ;
  END
END tt08-ssp-opamp
END LIBRARY

